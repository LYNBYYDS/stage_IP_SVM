----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 
-- Design Name: 
-- Module Name: TOP_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TOP_tb is
--  Port ( );
end TOP_tb;

architecture Behavioral of TOP_tb is

component TOP is 
	port (	-- SV
			SV0_dim0 : in std_logic_vector(27 downto 0); 
			SV0_dim1 : in std_logic_vector(27 downto 0); 
			SV0_dim2 : in std_logic_vector(27 downto 0); 
			SV0_dim3 : in std_logic_vector(27 downto 0); 
			SV0_dim4 : in std_logic_vector(27 downto 0); 
			SV0_dim5 : in std_logic_vector(27 downto 0); 
			SV0_dim6 : in std_logic_vector(27 downto 0); 
			SV0_dim7 : in std_logic_vector(27 downto 0); 
			SV1_dim0 : in std_logic_vector(27 downto 0); 
			SV1_dim1 : in std_logic_vector(27 downto 0); 
			SV1_dim2 : in std_logic_vector(27 downto 0); 
			SV1_dim3 : in std_logic_vector(27 downto 0); 
			SV1_dim4 : in std_logic_vector(27 downto 0); 
			SV1_dim5 : in std_logic_vector(27 downto 0); 
			SV1_dim6 : in std_logic_vector(27 downto 0); 
			SV1_dim7 : in std_logic_vector(27 downto 0); 
			SV2_dim0 : in std_logic_vector(27 downto 0); 
			SV2_dim1 : in std_logic_vector(27 downto 0); 
			SV2_dim2 : in std_logic_vector(27 downto 0); 
			SV2_dim3 : in std_logic_vector(27 downto 0); 
			SV2_dim4 : in std_logic_vector(27 downto 0); 
			SV2_dim5 : in std_logic_vector(27 downto 0); 
			SV2_dim6 : in std_logic_vector(27 downto 0); 
			SV2_dim7 : in std_logic_vector(27 downto 0); 
			SV3_dim0 : in std_logic_vector(27 downto 0); 
			SV3_dim1 : in std_logic_vector(27 downto 0); 
			SV3_dim2 : in std_logic_vector(27 downto 0); 
			SV3_dim3 : in std_logic_vector(27 downto 0); 
			SV3_dim4 : in std_logic_vector(27 downto 0); 
			SV3_dim5 : in std_logic_vector(27 downto 0); 
			SV3_dim6 : in std_logic_vector(27 downto 0); 
			SV3_dim7 : in std_logic_vector(27 downto 0); 
			SV4_dim0 : in std_logic_vector(27 downto 0); 
			SV4_dim1 : in std_logic_vector(27 downto 0); 
			SV4_dim2 : in std_logic_vector(27 downto 0); 
			SV4_dim3 : in std_logic_vector(27 downto 0); 
			SV4_dim4 : in std_logic_vector(27 downto 0); 
			SV4_dim5 : in std_logic_vector(27 downto 0); 
			SV4_dim6 : in std_logic_vector(27 downto 0); 
			SV4_dim7 : in std_logic_vector(27 downto 0); 
			SV5_dim0 : in std_logic_vector(27 downto 0); 
			SV5_dim1 : in std_logic_vector(27 downto 0); 
			SV5_dim2 : in std_logic_vector(27 downto 0); 
			SV5_dim3 : in std_logic_vector(27 downto 0); 
			SV5_dim4 : in std_logic_vector(27 downto 0); 
			SV5_dim5 : in std_logic_vector(27 downto 0); 
			SV5_dim6 : in std_logic_vector(27 downto 0); 
			SV5_dim7 : in std_logic_vector(27 downto 0); 
			SV6_dim0 : in std_logic_vector(27 downto 0); 
			SV6_dim1 : in std_logic_vector(27 downto 0); 
			SV6_dim2 : in std_logic_vector(27 downto 0); 
			SV6_dim3 : in std_logic_vector(27 downto 0); 
			SV6_dim4 : in std_logic_vector(27 downto 0); 
			SV6_dim5 : in std_logic_vector(27 downto 0); 
			SV6_dim6 : in std_logic_vector(27 downto 0); 
			SV6_dim7 : in std_logic_vector(27 downto 0); 
			SV7_dim0 : in std_logic_vector(27 downto 0); 
			SV7_dim1 : in std_logic_vector(27 downto 0); 
			SV7_dim2 : in std_logic_vector(27 downto 0); 
			SV7_dim3 : in std_logic_vector(27 downto 0); 
			SV7_dim4 : in std_logic_vector(27 downto 0); 
			SV7_dim5 : in std_logic_vector(27 downto 0); 
			SV7_dim6 : in std_logic_vector(27 downto 0); 
			SV7_dim7 : in std_logic_vector(27 downto 0); 
			SV8_dim0 : in std_logic_vector(27 downto 0); 
			SV8_dim1 : in std_logic_vector(27 downto 0); 
			SV8_dim2 : in std_logic_vector(27 downto 0); 
			SV8_dim3 : in std_logic_vector(27 downto 0); 
			SV8_dim4 : in std_logic_vector(27 downto 0); 
			SV8_dim5 : in std_logic_vector(27 downto 0); 
			SV8_dim6 : in std_logic_vector(27 downto 0); 
			SV8_dim7 : in std_logic_vector(27 downto 0); 
			SV9_dim0 : in std_logic_vector(27 downto 0); 
			SV9_dim1 : in std_logic_vector(27 downto 0); 
			SV9_dim2 : in std_logic_vector(27 downto 0); 
			SV9_dim3 : in std_logic_vector(27 downto 0); 
			SV9_dim4 : in std_logic_vector(27 downto 0); 
			SV9_dim5 : in std_logic_vector(27 downto 0); 
			SV9_dim6 : in std_logic_vector(27 downto 0); 
			SV9_dim7 : in std_logic_vector(27 downto 0); 
			SV10_dim0 : in std_logic_vector(27 downto 0); 
			SV10_dim1 : in std_logic_vector(27 downto 0); 
			SV10_dim2 : in std_logic_vector(27 downto 0); 
			SV10_dim3 : in std_logic_vector(27 downto 0); 
			SV10_dim4 : in std_logic_vector(27 downto 0); 
			SV10_dim5 : in std_logic_vector(27 downto 0); 
			SV10_dim6 : in std_logic_vector(27 downto 0); 
			SV10_dim7 : in std_logic_vector(27 downto 0); 
			SV11_dim0 : in std_logic_vector(27 downto 0); 
			SV11_dim1 : in std_logic_vector(27 downto 0); 
			SV11_dim2 : in std_logic_vector(27 downto 0); 
			SV11_dim3 : in std_logic_vector(27 downto 0); 
			SV11_dim4 : in std_logic_vector(27 downto 0); 
			SV11_dim5 : in std_logic_vector(27 downto 0); 
			SV11_dim6 : in std_logic_vector(27 downto 0); 
			SV11_dim7 : in std_logic_vector(27 downto 0); 
			SV12_dim0 : in std_logic_vector(27 downto 0); 
			SV12_dim1 : in std_logic_vector(27 downto 0); 
			SV12_dim2 : in std_logic_vector(27 downto 0); 
			SV12_dim3 : in std_logic_vector(27 downto 0); 
			SV12_dim4 : in std_logic_vector(27 downto 0); 
			SV12_dim5 : in std_logic_vector(27 downto 0); 
			SV12_dim6 : in std_logic_vector(27 downto 0); 
			SV12_dim7 : in std_logic_vector(27 downto 0); 
			SV13_dim0 : in std_logic_vector(27 downto 0); 
			SV13_dim1 : in std_logic_vector(27 downto 0); 
			SV13_dim2 : in std_logic_vector(27 downto 0); 
			SV13_dim3 : in std_logic_vector(27 downto 0); 
			SV13_dim4 : in std_logic_vector(27 downto 0); 
			SV13_dim5 : in std_logic_vector(27 downto 0); 
			SV13_dim6 : in std_logic_vector(27 downto 0); 
			SV13_dim7 : in std_logic_vector(27 downto 0); 
			SV14_dim0 : in std_logic_vector(27 downto 0); 
			SV14_dim1 : in std_logic_vector(27 downto 0); 
			SV14_dim2 : in std_logic_vector(27 downto 0); 
			SV14_dim3 : in std_logic_vector(27 downto 0); 
			SV14_dim4 : in std_logic_vector(27 downto 0); 
			SV14_dim5 : in std_logic_vector(27 downto 0); 
			SV14_dim6 : in std_logic_vector(27 downto 0); 
			SV14_dim7 : in std_logic_vector(27 downto 0); 
			SV15_dim0 : in std_logic_vector(27 downto 0); 
			SV15_dim1 : in std_logic_vector(27 downto 0); 
			SV15_dim2 : in std_logic_vector(27 downto 0); 
			SV15_dim3 : in std_logic_vector(27 downto 0); 
			SV15_dim4 : in std_logic_vector(27 downto 0); 
			SV15_dim5 : in std_logic_vector(27 downto 0); 
			SV15_dim6 : in std_logic_vector(27 downto 0); 
			SV15_dim7 : in std_logic_vector(27 downto 0); 
			SV16_dim0 : in std_logic_vector(27 downto 0); 
			SV16_dim1 : in std_logic_vector(27 downto 0); 
			SV16_dim2 : in std_logic_vector(27 downto 0); 
			SV16_dim3 : in std_logic_vector(27 downto 0); 
			SV16_dim4 : in std_logic_vector(27 downto 0); 
			SV16_dim5 : in std_logic_vector(27 downto 0); 
			SV16_dim6 : in std_logic_vector(27 downto 0); 
			SV16_dim7 : in std_logic_vector(27 downto 0); 
			SV17_dim0 : in std_logic_vector(27 downto 0); 
			SV17_dim1 : in std_logic_vector(27 downto 0); 
			SV17_dim2 : in std_logic_vector(27 downto 0); 
			SV17_dim3 : in std_logic_vector(27 downto 0); 
			SV17_dim4 : in std_logic_vector(27 downto 0); 
			SV17_dim5 : in std_logic_vector(27 downto 0); 
			SV17_dim6 : in std_logic_vector(27 downto 0); 
			SV17_dim7 : in std_logic_vector(27 downto 0); 
			SV18_dim0 : in std_logic_vector(27 downto 0); 
			SV18_dim1 : in std_logic_vector(27 downto 0); 
			SV18_dim2 : in std_logic_vector(27 downto 0); 
			SV18_dim3 : in std_logic_vector(27 downto 0); 
			SV18_dim4 : in std_logic_vector(27 downto 0); 
			SV18_dim5 : in std_logic_vector(27 downto 0); 
			SV18_dim6 : in std_logic_vector(27 downto 0); 
			SV18_dim7 : in std_logic_vector(27 downto 0); 
			SV19_dim0 : in std_logic_vector(27 downto 0); 
			SV19_dim1 : in std_logic_vector(27 downto 0); 
			SV19_dim2 : in std_logic_vector(27 downto 0); 
			SV19_dim3 : in std_logic_vector(27 downto 0); 
			SV19_dim4 : in std_logic_vector(27 downto 0); 
			SV19_dim5 : in std_logic_vector(27 downto 0); 
			SV19_dim6 : in std_logic_vector(27 downto 0); 
			SV19_dim7 : in std_logic_vector(27 downto 0); 
			SV20_dim0 : in std_logic_vector(27 downto 0); 
			SV20_dim1 : in std_logic_vector(27 downto 0); 
			SV20_dim2 : in std_logic_vector(27 downto 0); 
			SV20_dim3 : in std_logic_vector(27 downto 0); 
			SV20_dim4 : in std_logic_vector(27 downto 0); 
			SV20_dim5 : in std_logic_vector(27 downto 0); 
			SV20_dim6 : in std_logic_vector(27 downto 0); 
			SV20_dim7 : in std_logic_vector(27 downto 0); 
			SV21_dim0 : in std_logic_vector(27 downto 0); 
			SV21_dim1 : in std_logic_vector(27 downto 0); 
			SV21_dim2 : in std_logic_vector(27 downto 0); 
			SV21_dim3 : in std_logic_vector(27 downto 0); 
			SV21_dim4 : in std_logic_vector(27 downto 0); 
			SV21_dim5 : in std_logic_vector(27 downto 0); 
			SV21_dim6 : in std_logic_vector(27 downto 0); 
			SV21_dim7 : in std_logic_vector(27 downto 0); 
			SV22_dim0 : in std_logic_vector(27 downto 0); 
			SV22_dim1 : in std_logic_vector(27 downto 0); 
			SV22_dim2 : in std_logic_vector(27 downto 0); 
			SV22_dim3 : in std_logic_vector(27 downto 0); 
			SV22_dim4 : in std_logic_vector(27 downto 0); 
			SV22_dim5 : in std_logic_vector(27 downto 0); 
			SV22_dim6 : in std_logic_vector(27 downto 0); 
			SV22_dim7 : in std_logic_vector(27 downto 0); 
			SV23_dim0 : in std_logic_vector(27 downto 0); 
			SV23_dim1 : in std_logic_vector(27 downto 0); 
			SV23_dim2 : in std_logic_vector(27 downto 0); 
			SV23_dim3 : in std_logic_vector(27 downto 0); 
			SV23_dim4 : in std_logic_vector(27 downto 0); 
			SV23_dim5 : in std_logic_vector(27 downto 0); 
			SV23_dim6 : in std_logic_vector(27 downto 0); 
			SV23_dim7 : in std_logic_vector(27 downto 0); 
			SV24_dim0 : in std_logic_vector(27 downto 0); 
			SV24_dim1 : in std_logic_vector(27 downto 0); 
			SV24_dim2 : in std_logic_vector(27 downto 0); 
			SV24_dim3 : in std_logic_vector(27 downto 0); 
			SV24_dim4 : in std_logic_vector(27 downto 0); 
			SV24_dim5 : in std_logic_vector(27 downto 0); 
			SV24_dim6 : in std_logic_vector(27 downto 0); 
			SV24_dim7 : in std_logic_vector(27 downto 0); 
			SV25_dim0 : in std_logic_vector(27 downto 0); 
			SV25_dim1 : in std_logic_vector(27 downto 0); 
			SV25_dim2 : in std_logic_vector(27 downto 0); 
			SV25_dim3 : in std_logic_vector(27 downto 0); 
			SV25_dim4 : in std_logic_vector(27 downto 0); 
			SV25_dim5 : in std_logic_vector(27 downto 0); 
			SV25_dim6 : in std_logic_vector(27 downto 0); 
			SV25_dim7 : in std_logic_vector(27 downto 0); 
			SV26_dim0 : in std_logic_vector(27 downto 0); 
			SV26_dim1 : in std_logic_vector(27 downto 0); 
			SV26_dim2 : in std_logic_vector(27 downto 0); 
			SV26_dim3 : in std_logic_vector(27 downto 0); 
			SV26_dim4 : in std_logic_vector(27 downto 0); 
			SV26_dim5 : in std_logic_vector(27 downto 0); 
			SV26_dim6 : in std_logic_vector(27 downto 0); 
			SV26_dim7 : in std_logic_vector(27 downto 0); 
			SV27_dim0 : in std_logic_vector(27 downto 0); 
			SV27_dim1 : in std_logic_vector(27 downto 0); 
			SV27_dim2 : in std_logic_vector(27 downto 0); 
			SV27_dim3 : in std_logic_vector(27 downto 0); 
			SV27_dim4 : in std_logic_vector(27 downto 0); 
			SV27_dim5 : in std_logic_vector(27 downto 0); 
			SV27_dim6 : in std_logic_vector(27 downto 0); 
			SV27_dim7 : in std_logic_vector(27 downto 0); 
			SV28_dim0 : in std_logic_vector(27 downto 0); 
			SV28_dim1 : in std_logic_vector(27 downto 0); 
			SV28_dim2 : in std_logic_vector(27 downto 0); 
			SV28_dim3 : in std_logic_vector(27 downto 0); 
			SV28_dim4 : in std_logic_vector(27 downto 0); 
			SV28_dim5 : in std_logic_vector(27 downto 0); 
			SV28_dim6 : in std_logic_vector(27 downto 0); 
			SV28_dim7 : in std_logic_vector(27 downto 0); 
			SV29_dim0 : in std_logic_vector(27 downto 0); 
			SV29_dim1 : in std_logic_vector(27 downto 0); 
			SV29_dim2 : in std_logic_vector(27 downto 0); 
			SV29_dim3 : in std_logic_vector(27 downto 0); 
			SV29_dim4 : in std_logic_vector(27 downto 0); 
			SV29_dim5 : in std_logic_vector(27 downto 0); 
			SV29_dim6 : in std_logic_vector(27 downto 0); 
			SV29_dim7 : in std_logic_vector(27 downto 0); 
			SV30_dim0 : in std_logic_vector(27 downto 0); 
			SV30_dim1 : in std_logic_vector(27 downto 0); 
			SV30_dim2 : in std_logic_vector(27 downto 0); 
			SV30_dim3 : in std_logic_vector(27 downto 0); 
			SV30_dim4 : in std_logic_vector(27 downto 0); 
			SV30_dim5 : in std_logic_vector(27 downto 0); 
			SV30_dim6 : in std_logic_vector(27 downto 0); 
			SV30_dim7 : in std_logic_vector(27 downto 0); 
			SV31_dim0 : in std_logic_vector(27 downto 0); 
			SV31_dim1 : in std_logic_vector(27 downto 0); 
			SV31_dim2 : in std_logic_vector(27 downto 0); 
			SV31_dim3 : in std_logic_vector(27 downto 0); 
			SV31_dim4 : in std_logic_vector(27 downto 0); 
			SV31_dim5 : in std_logic_vector(27 downto 0); 
			SV31_dim6 : in std_logic_vector(27 downto 0); 
			SV31_dim7 : in std_logic_vector(27 downto 0); 
			SV32_dim0 : in std_logic_vector(27 downto 0); 
			SV32_dim1 : in std_logic_vector(27 downto 0); 
			SV32_dim2 : in std_logic_vector(27 downto 0); 
			SV32_dim3 : in std_logic_vector(27 downto 0); 
			SV32_dim4 : in std_logic_vector(27 downto 0); 
			SV32_dim5 : in std_logic_vector(27 downto 0); 
			SV32_dim6 : in std_logic_vector(27 downto 0); 
			SV32_dim7 : in std_logic_vector(27 downto 0); 
			SV33_dim0 : in std_logic_vector(27 downto 0); 
			SV33_dim1 : in std_logic_vector(27 downto 0); 
			SV33_dim2 : in std_logic_vector(27 downto 0); 
			SV33_dim3 : in std_logic_vector(27 downto 0); 
			SV33_dim4 : in std_logic_vector(27 downto 0); 
			SV33_dim5 : in std_logic_vector(27 downto 0); 
			SV33_dim6 : in std_logic_vector(27 downto 0); 
			SV33_dim7 : in std_logic_vector(27 downto 0); 
			SV34_dim0 : in std_logic_vector(27 downto 0); 
			SV34_dim1 : in std_logic_vector(27 downto 0); 
			SV34_dim2 : in std_logic_vector(27 downto 0); 
			SV34_dim3 : in std_logic_vector(27 downto 0); 
			SV34_dim4 : in std_logic_vector(27 downto 0); 
			SV34_dim5 : in std_logic_vector(27 downto 0); 
			SV34_dim6 : in std_logic_vector(27 downto 0); 
			SV34_dim7 : in std_logic_vector(27 downto 0); 
			SV35_dim0 : in std_logic_vector(27 downto 0); 
			SV35_dim1 : in std_logic_vector(27 downto 0); 
			SV35_dim2 : in std_logic_vector(27 downto 0); 
			SV35_dim3 : in std_logic_vector(27 downto 0); 
			SV35_dim4 : in std_logic_vector(27 downto 0); 
			SV35_dim5 : in std_logic_vector(27 downto 0); 
			SV35_dim6 : in std_logic_vector(27 downto 0); 
			SV35_dim7 : in std_logic_vector(27 downto 0); 
			SV36_dim0 : in std_logic_vector(27 downto 0); 
			SV36_dim1 : in std_logic_vector(27 downto 0); 
			SV36_dim2 : in std_logic_vector(27 downto 0); 
			SV36_dim3 : in std_logic_vector(27 downto 0); 
			SV36_dim4 : in std_logic_vector(27 downto 0); 
			SV36_dim5 : in std_logic_vector(27 downto 0); 
			SV36_dim6 : in std_logic_vector(27 downto 0); 
			SV36_dim7 : in std_logic_vector(27 downto 0); 
			SV37_dim0 : in std_logic_vector(27 downto 0); 
			SV37_dim1 : in std_logic_vector(27 downto 0); 
			SV37_dim2 : in std_logic_vector(27 downto 0); 
			SV37_dim3 : in std_logic_vector(27 downto 0); 
			SV37_dim4 : in std_logic_vector(27 downto 0); 
			SV37_dim5 : in std_logic_vector(27 downto 0); 
			SV37_dim6 : in std_logic_vector(27 downto 0); 
			SV37_dim7 : in std_logic_vector(27 downto 0); 
			SV38_dim0 : in std_logic_vector(27 downto 0); 
			SV38_dim1 : in std_logic_vector(27 downto 0); 
			SV38_dim2 : in std_logic_vector(27 downto 0); 
			SV38_dim3 : in std_logic_vector(27 downto 0); 
			SV38_dim4 : in std_logic_vector(27 downto 0); 
			SV38_dim5 : in std_logic_vector(27 downto 0); 
			SV38_dim6 : in std_logic_vector(27 downto 0); 
			SV38_dim7 : in std_logic_vector(27 downto 0); 
			SV39_dim0 : in std_logic_vector(27 downto 0); 
			SV39_dim1 : in std_logic_vector(27 downto 0); 
			SV39_dim2 : in std_logic_vector(27 downto 0); 
			SV39_dim3 : in std_logic_vector(27 downto 0); 
			SV39_dim4 : in std_logic_vector(27 downto 0); 
			SV39_dim5 : in std_logic_vector(27 downto 0); 
			SV39_dim6 : in std_logic_vector(27 downto 0); 
			SV39_dim7 : in std_logic_vector(27 downto 0); 
			SV40_dim0 : in std_logic_vector(27 downto 0); 
			SV40_dim1 : in std_logic_vector(27 downto 0); 
			SV40_dim2 : in std_logic_vector(27 downto 0); 
			SV40_dim3 : in std_logic_vector(27 downto 0); 
			SV40_dim4 : in std_logic_vector(27 downto 0); 
			SV40_dim5 : in std_logic_vector(27 downto 0); 
			SV40_dim6 : in std_logic_vector(27 downto 0); 
			SV40_dim7 : in std_logic_vector(27 downto 0); 
			SV41_dim0 : in std_logic_vector(27 downto 0); 
			SV41_dim1 : in std_logic_vector(27 downto 0); 
			SV41_dim2 : in std_logic_vector(27 downto 0); 
			SV41_dim3 : in std_logic_vector(27 downto 0); 
			SV41_dim4 : in std_logic_vector(27 downto 0); 
			SV41_dim5 : in std_logic_vector(27 downto 0); 
			SV41_dim6 : in std_logic_vector(27 downto 0); 
			SV41_dim7 : in std_logic_vector(27 downto 0); 
			SV42_dim0 : in std_logic_vector(27 downto 0); 
			SV42_dim1 : in std_logic_vector(27 downto 0); 
			SV42_dim2 : in std_logic_vector(27 downto 0); 
			SV42_dim3 : in std_logic_vector(27 downto 0); 
			SV42_dim4 : in std_logic_vector(27 downto 0); 
			SV42_dim5 : in std_logic_vector(27 downto 0); 
			SV42_dim6 : in std_logic_vector(27 downto 0); 
			SV42_dim7 : in std_logic_vector(27 downto 0); 
			SV43_dim0 : in std_logic_vector(27 downto 0); 
			SV43_dim1 : in std_logic_vector(27 downto 0); 
			SV43_dim2 : in std_logic_vector(27 downto 0); 
			SV43_dim3 : in std_logic_vector(27 downto 0); 
			SV43_dim4 : in std_logic_vector(27 downto 0); 
			SV43_dim5 : in std_logic_vector(27 downto 0); 
			SV43_dim6 : in std_logic_vector(27 downto 0); 
			SV43_dim7 : in std_logic_vector(27 downto 0); 
			SV44_dim0 : in std_logic_vector(27 downto 0); 
			SV44_dim1 : in std_logic_vector(27 downto 0); 
			SV44_dim2 : in std_logic_vector(27 downto 0); 
			SV44_dim3 : in std_logic_vector(27 downto 0); 
			SV44_dim4 : in std_logic_vector(27 downto 0); 
			SV44_dim5 : in std_logic_vector(27 downto 0); 
			SV44_dim6 : in std_logic_vector(27 downto 0); 
			SV44_dim7 : in std_logic_vector(27 downto 0); 
			SV45_dim0 : in std_logic_vector(27 downto 0); 
			SV45_dim1 : in std_logic_vector(27 downto 0); 
			SV45_dim2 : in std_logic_vector(27 downto 0); 
			SV45_dim3 : in std_logic_vector(27 downto 0); 
			SV45_dim4 : in std_logic_vector(27 downto 0); 
			SV45_dim5 : in std_logic_vector(27 downto 0); 
			SV45_dim6 : in std_logic_vector(27 downto 0); 
			SV45_dim7 : in std_logic_vector(27 downto 0); 
			SV46_dim0 : in std_logic_vector(27 downto 0); 
			SV46_dim1 : in std_logic_vector(27 downto 0); 
			SV46_dim2 : in std_logic_vector(27 downto 0); 
			SV46_dim3 : in std_logic_vector(27 downto 0); 
			SV46_dim4 : in std_logic_vector(27 downto 0); 
			SV46_dim5 : in std_logic_vector(27 downto 0); 
			SV46_dim6 : in std_logic_vector(27 downto 0); 
			SV46_dim7 : in std_logic_vector(27 downto 0); 
			SV47_dim0 : in std_logic_vector(27 downto 0); 
			SV47_dim1 : in std_logic_vector(27 downto 0); 
			SV47_dim2 : in std_logic_vector(27 downto 0); 
			SV47_dim3 : in std_logic_vector(27 downto 0); 
			SV47_dim4 : in std_logic_vector(27 downto 0); 
			SV47_dim5 : in std_logic_vector(27 downto 0); 
			SV47_dim6 : in std_logic_vector(27 downto 0); 
			SV47_dim7 : in std_logic_vector(27 downto 0); 
			SV48_dim0 : in std_logic_vector(27 downto 0); 
			SV48_dim1 : in std_logic_vector(27 downto 0); 
			SV48_dim2 : in std_logic_vector(27 downto 0); 
			SV48_dim3 : in std_logic_vector(27 downto 0); 
			SV48_dim4 : in std_logic_vector(27 downto 0); 
			SV48_dim5 : in std_logic_vector(27 downto 0); 
			SV48_dim6 : in std_logic_vector(27 downto 0); 
			SV48_dim7 : in std_logic_vector(27 downto 0); 
			SV49_dim0 : in std_logic_vector(27 downto 0); 
			SV49_dim1 : in std_logic_vector(27 downto 0); 
			SV49_dim2 : in std_logic_vector(27 downto 0); 
			SV49_dim3 : in std_logic_vector(27 downto 0); 
			SV49_dim4 : in std_logic_vector(27 downto 0); 
			SV49_dim5 : in std_logic_vector(27 downto 0); 
			SV49_dim6 : in std_logic_vector(27 downto 0); 
			SV49_dim7 : in std_logic_vector(27 downto 0); 
			SV50_dim0 : in std_logic_vector(27 downto 0); 
			SV50_dim1 : in std_logic_vector(27 downto 0); 
			SV50_dim2 : in std_logic_vector(27 downto 0); 
			SV50_dim3 : in std_logic_vector(27 downto 0); 
			SV50_dim4 : in std_logic_vector(27 downto 0); 
			SV50_dim5 : in std_logic_vector(27 downto 0); 
			SV50_dim6 : in std_logic_vector(27 downto 0); 
			SV50_dim7 : in std_logic_vector(27 downto 0); 
			SV51_dim0 : in std_logic_vector(27 downto 0); 
			SV51_dim1 : in std_logic_vector(27 downto 0); 
			SV51_dim2 : in std_logic_vector(27 downto 0); 
			SV51_dim3 : in std_logic_vector(27 downto 0); 
			SV51_dim4 : in std_logic_vector(27 downto 0); 
			SV51_dim5 : in std_logic_vector(27 downto 0); 
			SV51_dim6 : in std_logic_vector(27 downto 0); 
			SV51_dim7 : in std_logic_vector(27 downto 0); 
			SV52_dim0 : in std_logic_vector(27 downto 0); 
			SV52_dim1 : in std_logic_vector(27 downto 0); 
			SV52_dim2 : in std_logic_vector(27 downto 0); 
			SV52_dim3 : in std_logic_vector(27 downto 0); 
			SV52_dim4 : in std_logic_vector(27 downto 0); 
			SV52_dim5 : in std_logic_vector(27 downto 0); 
			SV52_dim6 : in std_logic_vector(27 downto 0); 
			SV52_dim7 : in std_logic_vector(27 downto 0); 
			SV53_dim0 : in std_logic_vector(27 downto 0); 
			SV53_dim1 : in std_logic_vector(27 downto 0); 
			SV53_dim2 : in std_logic_vector(27 downto 0); 
			SV53_dim3 : in std_logic_vector(27 downto 0); 
			SV53_dim4 : in std_logic_vector(27 downto 0); 
			SV53_dim5 : in std_logic_vector(27 downto 0); 
			SV53_dim6 : in std_logic_vector(27 downto 0); 
			SV53_dim7 : in std_logic_vector(27 downto 0); 
			SV54_dim0 : in std_logic_vector(27 downto 0); 
			SV54_dim1 : in std_logic_vector(27 downto 0); 
			SV54_dim2 : in std_logic_vector(27 downto 0); 
			SV54_dim3 : in std_logic_vector(27 downto 0); 
			SV54_dim4 : in std_logic_vector(27 downto 0); 
			SV54_dim5 : in std_logic_vector(27 downto 0); 
			SV54_dim6 : in std_logic_vector(27 downto 0); 
			SV54_dim7 : in std_logic_vector(27 downto 0); 
			SV55_dim0 : in std_logic_vector(27 downto 0); 
			SV55_dim1 : in std_logic_vector(27 downto 0); 
			SV55_dim2 : in std_logic_vector(27 downto 0); 
			SV55_dim3 : in std_logic_vector(27 downto 0); 
			SV55_dim4 : in std_logic_vector(27 downto 0); 
			SV55_dim5 : in std_logic_vector(27 downto 0); 
			SV55_dim6 : in std_logic_vector(27 downto 0); 
			SV55_dim7 : in std_logic_vector(27 downto 0); 
			SV56_dim0 : in std_logic_vector(27 downto 0); 
			SV56_dim1 : in std_logic_vector(27 downto 0); 
			SV56_dim2 : in std_logic_vector(27 downto 0); 
			SV56_dim3 : in std_logic_vector(27 downto 0); 
			SV56_dim4 : in std_logic_vector(27 downto 0); 
			SV56_dim5 : in std_logic_vector(27 downto 0); 
			SV56_dim6 : in std_logic_vector(27 downto 0); 
			SV56_dim7 : in std_logic_vector(27 downto 0); 
			SV57_dim0 : in std_logic_vector(27 downto 0); 
			SV57_dim1 : in std_logic_vector(27 downto 0); 
			SV57_dim2 : in std_logic_vector(27 downto 0); 
			SV57_dim3 : in std_logic_vector(27 downto 0); 
			SV57_dim4 : in std_logic_vector(27 downto 0); 
			SV57_dim5 : in std_logic_vector(27 downto 0); 
			SV57_dim6 : in std_logic_vector(27 downto 0); 
			SV57_dim7 : in std_logic_vector(27 downto 0); 
			SV58_dim0 : in std_logic_vector(27 downto 0); 
			SV58_dim1 : in std_logic_vector(27 downto 0); 
			SV58_dim2 : in std_logic_vector(27 downto 0); 
			SV58_dim3 : in std_logic_vector(27 downto 0); 
			SV58_dim4 : in std_logic_vector(27 downto 0); 
			SV58_dim5 : in std_logic_vector(27 downto 0); 
			SV58_dim6 : in std_logic_vector(27 downto 0); 
			SV58_dim7 : in std_logic_vector(27 downto 0); 
			SV59_dim0 : in std_logic_vector(27 downto 0); 
			SV59_dim1 : in std_logic_vector(27 downto 0); 
			SV59_dim2 : in std_logic_vector(27 downto 0); 
			SV59_dim3 : in std_logic_vector(27 downto 0); 
			SV59_dim4 : in std_logic_vector(27 downto 0); 
			SV59_dim5 : in std_logic_vector(27 downto 0); 
			SV59_dim6 : in std_logic_vector(27 downto 0); 
			SV59_dim7 : in std_logic_vector(27 downto 0); 
			SV60_dim0 : in std_logic_vector(27 downto 0); 
			SV60_dim1 : in std_logic_vector(27 downto 0); 
			SV60_dim2 : in std_logic_vector(27 downto 0); 
			SV60_dim3 : in std_logic_vector(27 downto 0); 
			SV60_dim4 : in std_logic_vector(27 downto 0); 
			SV60_dim5 : in std_logic_vector(27 downto 0); 
			SV60_dim6 : in std_logic_vector(27 downto 0); 
			SV60_dim7 : in std_logic_vector(27 downto 0); 
			SV61_dim0 : in std_logic_vector(27 downto 0); 
			SV61_dim1 : in std_logic_vector(27 downto 0); 
			SV61_dim2 : in std_logic_vector(27 downto 0); 
			SV61_dim3 : in std_logic_vector(27 downto 0); 
			SV61_dim4 : in std_logic_vector(27 downto 0); 
			SV61_dim5 : in std_logic_vector(27 downto 0); 
			SV61_dim6 : in std_logic_vector(27 downto 0); 
			SV61_dim7 : in std_logic_vector(27 downto 0); 
			SV62_dim0 : in std_logic_vector(27 downto 0); 
			SV62_dim1 : in std_logic_vector(27 downto 0); 
			SV62_dim2 : in std_logic_vector(27 downto 0); 
			SV62_dim3 : in std_logic_vector(27 downto 0); 
			SV62_dim4 : in std_logic_vector(27 downto 0); 
			SV62_dim5 : in std_logic_vector(27 downto 0); 
			SV62_dim6 : in std_logic_vector(27 downto 0); 
			SV62_dim7 : in std_logic_vector(27 downto 0); 
			SV63_dim0 : in std_logic_vector(27 downto 0); 
			SV63_dim1 : in std_logic_vector(27 downto 0); 
			SV63_dim2 : in std_logic_vector(27 downto 0); 
			SV63_dim3 : in std_logic_vector(27 downto 0); 
			SV63_dim4 : in std_logic_vector(27 downto 0); 
			SV63_dim5 : in std_logic_vector(27 downto 0); 
			SV63_dim6 : in std_logic_vector(27 downto 0); 
			SV63_dim7 : in std_logic_vector(27 downto 0); 
			SV64_dim0 : in std_logic_vector(27 downto 0); 
			SV64_dim1 : in std_logic_vector(27 downto 0); 
			SV64_dim2 : in std_logic_vector(27 downto 0); 
			SV64_dim3 : in std_logic_vector(27 downto 0); 
			SV64_dim4 : in std_logic_vector(27 downto 0); 
			SV64_dim5 : in std_logic_vector(27 downto 0); 
			SV64_dim6 : in std_logic_vector(27 downto 0); 
			SV64_dim7 : in std_logic_vector(27 downto 0); 
			SV65_dim0 : in std_logic_vector(27 downto 0); 
			SV65_dim1 : in std_logic_vector(27 downto 0); 
			SV65_dim2 : in std_logic_vector(27 downto 0); 
			SV65_dim3 : in std_logic_vector(27 downto 0); 
			SV65_dim4 : in std_logic_vector(27 downto 0); 
			SV65_dim5 : in std_logic_vector(27 downto 0); 
			SV65_dim6 : in std_logic_vector(27 downto 0); 
			SV65_dim7 : in std_logic_vector(27 downto 0); 
			SV66_dim0 : in std_logic_vector(27 downto 0); 
			SV66_dim1 : in std_logic_vector(27 downto 0); 
			SV66_dim2 : in std_logic_vector(27 downto 0); 
			SV66_dim3 : in std_logic_vector(27 downto 0); 
			SV66_dim4 : in std_logic_vector(27 downto 0); 
			SV66_dim5 : in std_logic_vector(27 downto 0); 
			SV66_dim6 : in std_logic_vector(27 downto 0); 
			SV66_dim7 : in std_logic_vector(27 downto 0); 
			SV67_dim0 : in std_logic_vector(27 downto 0); 
			SV67_dim1 : in std_logic_vector(27 downto 0); 
			SV67_dim2 : in std_logic_vector(27 downto 0); 
			SV67_dim3 : in std_logic_vector(27 downto 0); 
			SV67_dim4 : in std_logic_vector(27 downto 0); 
			SV67_dim5 : in std_logic_vector(27 downto 0); 
			SV67_dim6 : in std_logic_vector(27 downto 0); 
			SV67_dim7 : in std_logic_vector(27 downto 0); 
			SV68_dim0 : in std_logic_vector(27 downto 0); 
			SV68_dim1 : in std_logic_vector(27 downto 0); 
			SV68_dim2 : in std_logic_vector(27 downto 0); 
			SV68_dim3 : in std_logic_vector(27 downto 0); 
			SV68_dim4 : in std_logic_vector(27 downto 0); 
			SV68_dim5 : in std_logic_vector(27 downto 0); 
			SV68_dim6 : in std_logic_vector(27 downto 0); 
			SV68_dim7 : in std_logic_vector(27 downto 0); 
			SV69_dim0 : in std_logic_vector(27 downto 0); 
			SV69_dim1 : in std_logic_vector(27 downto 0); 
			SV69_dim2 : in std_logic_vector(27 downto 0); 
			SV69_dim3 : in std_logic_vector(27 downto 0); 
			SV69_dim4 : in std_logic_vector(27 downto 0); 
			SV69_dim5 : in std_logic_vector(27 downto 0); 
			SV69_dim6 : in std_logic_vector(27 downto 0); 
			SV69_dim7 : in std_logic_vector(27 downto 0); 
			SV70_dim0 : in std_logic_vector(27 downto 0); 
			SV70_dim1 : in std_logic_vector(27 downto 0); 
			SV70_dim2 : in std_logic_vector(27 downto 0); 
			SV70_dim3 : in std_logic_vector(27 downto 0); 
			SV70_dim4 : in std_logic_vector(27 downto 0); 
			SV70_dim5 : in std_logic_vector(27 downto 0); 
			SV70_dim6 : in std_logic_vector(27 downto 0); 
			SV70_dim7 : in std_logic_vector(27 downto 0); 

			-- Test Data
			test_data_dim0 : in std_logic_vector(27 downto 0); 
			test_data_dim1 : in std_logic_vector(27 downto 0); 
			test_data_dim2 : in std_logic_vector(27 downto 0); 
			test_data_dim3 : in std_logic_vector(27 downto 0); 
			test_data_dim4 : in std_logic_vector(27 downto 0); 
			test_data_dim5 : in std_logic_vector(27 downto 0); 
			test_data_dim6 : in std_logic_vector(27 downto 0); 
			test_data_dim7 : in std_logic_vector(27 downto 0); 

			-- alpha * Y
			SV0_alphaY : in std_logic_vector(11 downto 0); 
			SV1_alphaY : in std_logic_vector(11 downto 0); 
			SV2_alphaY : in std_logic_vector(11 downto 0); 
			SV3_alphaY : in std_logic_vector(11 downto 0); 
			SV4_alphaY : in std_logic_vector(11 downto 0); 
			SV5_alphaY : in std_logic_vector(11 downto 0); 
			SV6_alphaY : in std_logic_vector(11 downto 0); 
			SV7_alphaY : in std_logic_vector(11 downto 0); 
			SV8_alphaY : in std_logic_vector(11 downto 0); 
			SV9_alphaY : in std_logic_vector(11 downto 0); 
			SV10_alphaY : in std_logic_vector(11 downto 0); 
			SV11_alphaY : in std_logic_vector(11 downto 0); 
			SV12_alphaY : in std_logic_vector(11 downto 0); 
			SV13_alphaY : in std_logic_vector(11 downto 0); 
			SV14_alphaY : in std_logic_vector(11 downto 0); 
			SV15_alphaY : in std_logic_vector(11 downto 0); 
			SV16_alphaY : in std_logic_vector(11 downto 0); 
			SV17_alphaY : in std_logic_vector(11 downto 0); 
			SV18_alphaY : in std_logic_vector(11 downto 0); 
			SV19_alphaY : in std_logic_vector(11 downto 0); 
			SV20_alphaY : in std_logic_vector(11 downto 0); 
			SV21_alphaY : in std_logic_vector(11 downto 0); 
			SV22_alphaY : in std_logic_vector(11 downto 0); 
			SV23_alphaY : in std_logic_vector(11 downto 0); 
			SV24_alphaY : in std_logic_vector(11 downto 0); 
			SV25_alphaY : in std_logic_vector(11 downto 0); 
			SV26_alphaY : in std_logic_vector(11 downto 0); 
			SV27_alphaY : in std_logic_vector(11 downto 0); 
			SV28_alphaY : in std_logic_vector(11 downto 0); 
			SV29_alphaY : in std_logic_vector(11 downto 0); 
			SV30_alphaY : in std_logic_vector(11 downto 0); 
			SV31_alphaY : in std_logic_vector(11 downto 0); 
			SV32_alphaY : in std_logic_vector(11 downto 0); 
			SV33_alphaY : in std_logic_vector(11 downto 0); 
			SV34_alphaY : in std_logic_vector(11 downto 0); 
			SV35_alphaY : in std_logic_vector(11 downto 0); 
			SV36_alphaY : in std_logic_vector(11 downto 0); 
			SV37_alphaY : in std_logic_vector(11 downto 0); 
			SV38_alphaY : in std_logic_vector(11 downto 0); 
			SV39_alphaY : in std_logic_vector(11 downto 0); 
			SV40_alphaY : in std_logic_vector(11 downto 0); 
			SV41_alphaY : in std_logic_vector(11 downto 0); 
			SV42_alphaY : in std_logic_vector(11 downto 0); 
			SV43_alphaY : in std_logic_vector(11 downto 0); 
			SV44_alphaY : in std_logic_vector(11 downto 0); 
			SV45_alphaY : in std_logic_vector(11 downto 0); 
			SV46_alphaY : in std_logic_vector(11 downto 0); 
			SV47_alphaY : in std_logic_vector(11 downto 0); 
			SV48_alphaY : in std_logic_vector(11 downto 0); 
			SV49_alphaY : in std_logic_vector(11 downto 0); 
			SV50_alphaY : in std_logic_vector(11 downto 0); 
			SV51_alphaY : in std_logic_vector(11 downto 0); 
			SV52_alphaY : in std_logic_vector(11 downto 0); 
			SV53_alphaY : in std_logic_vector(11 downto 0); 
			SV54_alphaY : in std_logic_vector(11 downto 0); 
			SV55_alphaY : in std_logic_vector(11 downto 0); 
			SV56_alphaY : in std_logic_vector(11 downto 0); 
			SV57_alphaY : in std_logic_vector(11 downto 0); 
			SV58_alphaY : in std_logic_vector(11 downto 0); 
			SV59_alphaY : in std_logic_vector(11 downto 0); 
			SV60_alphaY : in std_logic_vector(11 downto 0); 
			SV61_alphaY : in std_logic_vector(11 downto 0); 
			SV62_alphaY : in std_logic_vector(11 downto 0); 
			SV63_alphaY : in std_logic_vector(11 downto 0); 
			SV64_alphaY : in std_logic_vector(11 downto 0); 
			SV65_alphaY : in std_logic_vector(11 downto 0); 
			SV66_alphaY : in std_logic_vector(11 downto 0); 
			SV67_alphaY : in std_logic_vector(11 downto 0); 
			SV68_alphaY : in std_logic_vector(11 downto 0); 
			SV69_alphaY : in std_logic_vector(11 downto 0); 
			SV70_alphaY : in std_logic_vector(11 downto 0); 

			-- gamma
			gamma : in std_logic_vector(11 downto 0); 

			-- b
			b : in std_logic_vector(19 downto 0); 

			-- output
			output : out std_logic 
			);
end component;

signal SV0_dim0 : std_logic_vector(27 downto 0) := "0001100100010100110110111000";
signal SV0_dim1 : std_logic_vector(27 downto 0) := "0000000000000111110100010100";
signal SV0_dim2 : std_logic_vector(27 downto 0) := "0000000011001101010101010010";
signal SV0_dim3 : std_logic_vector(27 downto 0) := "0000000010010010001100010100";
signal SV0_dim4 : std_logic_vector(27 downto 0) := "0000000000110010101100011111";
signal SV0_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110101010010";
signal SV0_dim6 : std_logic_vector(27 downto 0) := "0000000000000000010111001101";
signal SV0_dim7 : std_logic_vector(27 downto 0) := "0000000000001010010000111101";
signal SV1_dim0 : std_logic_vector(27 downto 0) := "0001101000011010110001100110";
signal SV1_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100100101001";
signal SV1_dim2 : std_logic_vector(27 downto 0) := "0000000010000100111000111101";
signal SV1_dim3 : std_logic_vector(27 downto 0) := "0000000010000000010100110011";
signal SV1_dim4 : std_logic_vector(27 downto 0) := "0000000111110001100110111000";
signal SV1_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV1_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV1_dim7 : std_logic_vector(27 downto 0) := "0000000000000010111000001010";
signal SV2_dim0 : std_logic_vector(27 downto 0) := "0010000111110111000001011100";
signal SV2_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101001100110";
signal SV2_dim2 : std_logic_vector(27 downto 0) := "0000000100011100001010101110";
signal SV2_dim3 : std_logic_vector(27 downto 0) := "0000000010010000100111010111";
signal SV2_dim4 : std_logic_vector(27 downto 0) := "0000000000101110000111100001";
signal SV2_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110000110011";
signal SV2_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110011010";
signal SV2_dim7 : std_logic_vector(27 downto 0) := "0000000000001010101001011100";
signal SV3_dim0 : std_logic_vector(27 downto 0) := "0010101110010110110111001101";
signal SV3_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101011100001";
signal SV3_dim2 : std_logic_vector(27 downto 0) := "0000000011011100000000000000";
signal SV3_dim3 : std_logic_vector(27 downto 0) := "0000000010000101010100010100";
signal SV3_dim4 : std_logic_vector(27 downto 0) := "0000000111110010001010001111";
signal SV3_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV3_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV3_dim7 : std_logic_vector(27 downto 0) := "0000000000000010111111001101";
signal SV4_dim0 : std_logic_vector(27 downto 0) := "0001010001010001101101110001";
signal SV4_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101001100110";
signal SV4_dim2 : std_logic_vector(27 downto 0) := "0000000010101010000000000000";
signal SV4_dim3 : std_logic_vector(27 downto 0) := "0000000010010011100111110110";
signal SV4_dim4 : std_logic_vector(27 downto 0) := "0000000000110001000110111000";
signal SV4_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110011100001";
signal SV4_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011001110001";
signal SV4_dim7 : std_logic_vector(27 downto 0) := "0000000000001010100010000101";
signal SV5_dim0 : std_logic_vector(27 downto 0) := "0001100110110110001100101001";
signal SV5_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100100101001";
signal SV5_dim2 : std_logic_vector(27 downto 0) := "0000000010000010111000111101";
signal SV5_dim3 : std_logic_vector(27 downto 0) := "0000000010000101000100110011";
signal SV5_dim4 : std_logic_vector(27 downto 0) := "0000000111110001100110111000";
signal SV5_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV5_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV5_dim7 : std_logic_vector(27 downto 0) := "0000000000000010111110111000";
signal SV6_dim0 : std_logic_vector(27 downto 0) := "0010110000101011001000000000";
signal SV6_dim1 : std_logic_vector(27 downto 0) := "0000000000001010000110000101";
signal SV6_dim2 : std_logic_vector(27 downto 0) := "0000000100011000000000000000";
signal SV6_dim3 : std_logic_vector(27 downto 0) := "0000000010010000100011101100";
signal SV6_dim4 : std_logic_vector(27 downto 0) := "0000000100100001000101001000";
signal SV6_dim5 : std_logic_vector(27 downto 0) := "0000000000000000001011110110";
signal SV6_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011010101110";
signal SV6_dim7 : std_logic_vector(27 downto 0) := "0000000000000100010000000000";
signal SV7_dim0 : std_logic_vector(27 downto 0) := "0010101001110101010100101001";
signal SV7_dim1 : std_logic_vector(27 downto 0) := "0000000000000111111000001010";
signal SV7_dim2 : std_logic_vector(27 downto 0) := "0000000101011001000000000000";
signal SV7_dim3 : std_logic_vector(27 downto 0) := "0000000001110011000011100001";
signal SV7_dim4 : std_logic_vector(27 downto 0) := "0000000010101110011001011100";
signal SV7_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100101001";
signal SV7_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101010101110";
signal SV7_dim7 : std_logic_vector(27 downto 0) := "0000000000000100010110101110";
signal SV8_dim0 : std_logic_vector(27 downto 0) := "0001010100110010010001100110";
signal SV8_dim1 : std_logic_vector(27 downto 0) := "0000000000001010001100110011";
signal SV8_dim2 : std_logic_vector(27 downto 0) := "0000000010000101000000000000";
signal SV8_dim3 : std_logic_vector(27 downto 0) := "0000000001110001010101100110";
signal SV8_dim4 : std_logic_vector(27 downto 0) := "0000000001011010100010100100";
signal SV8_dim5 : std_logic_vector(27 downto 0) := "0000000000000000001011010111";
signal SV8_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011000000000";
signal SV8_dim7 : std_logic_vector(27 downto 0) := "0000000000000101111101001000";
signal SV9_dim0 : std_logic_vector(27 downto 0) := "0000001110111000111111110110";
signal SV9_dim1 : std_logic_vector(27 downto 0) := "0000000000000011110010111000";
signal SV9_dim2 : std_logic_vector(27 downto 0) := "0000000000111110110010111000";
signal SV9_dim3 : std_logic_vector(27 downto 0) := "0000000001101110010000101001";
signal SV9_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000001010010";
signal SV9_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111111001101";
signal SV9_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110001111";
signal SV9_dim7 : std_logic_vector(27 downto 0) := "0000000110000001000000011111";
signal SV10_dim0 : std_logic_vector(27 downto 0) := "0001001110011000101010101110";
signal SV10_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV10_dim2 : std_logic_vector(27 downto 0) := "0000000001100100010101010010";
signal SV10_dim3 : std_logic_vector(27 downto 0) := "0000000010000011011011010111";
signal SV10_dim4 : std_logic_vector(27 downto 0) := "0000000001101011001001001000";
signal SV10_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010110001111";
signal SV10_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101111000011";
signal SV10_dim7 : std_logic_vector(27 downto 0) := "0000000000000110010110001111";
signal SV11_dim0 : std_logic_vector(27 downto 0) := "0001001111110101010100000000";
signal SV11_dim1 : std_logic_vector(27 downto 0) := "0000000000000111110000011111";
signal SV11_dim2 : std_logic_vector(27 downto 0) := "0000000010100100101010101110";
signal SV11_dim3 : std_logic_vector(27 downto 0) := "0000000010010101001000010100";
signal SV11_dim4 : std_logic_vector(27 downto 0) := "0000000000110000110000111101";
signal SV11_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110011010111";
signal SV11_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011010000101";
signal SV11_dim7 : std_logic_vector(27 downto 0) := "0000000000001010101011010111";
signal SV12_dim0 : std_logic_vector(27 downto 0) := "0001011100111110000000000000";
signal SV12_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV12_dim2 : std_logic_vector(27 downto 0) := "0000000001110111000000000000";
signal SV12_dim3 : std_logic_vector(27 downto 0) := "0000000010001110010001001000";
signal SV12_dim4 : std_logic_vector(27 downto 0) := "0000000001110100011101001000";
signal SV12_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010011010111";
signal SV12_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111010111";
signal SV12_dim7 : std_logic_vector(27 downto 0) := "0000000000000110100101111011";
signal SV13_dim0 : std_logic_vector(27 downto 0) := "0001101100011011110011100001";
signal SV13_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100100101001";
signal SV13_dim2 : std_logic_vector(27 downto 0) := "0000000010001010000000000000";
signal SV13_dim3 : std_logic_vector(27 downto 0) := "0000000001111001000100110011";
signal SV13_dim4 : std_logic_vector(27 downto 0) := "0000000111110001100110111000";
signal SV13_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV13_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV13_dim7 : std_logic_vector(27 downto 0) := "0000000000000010101101110001";
signal SV14_dim0 : std_logic_vector(27 downto 0) := "0010000110001000110100010100";
signal SV14_dim1 : std_logic_vector(27 downto 0) := "0000000000000011111011101100";
signal SV14_dim2 : std_logic_vector(27 downto 0) := "0000001000100001110110111000";
signal SV14_dim3 : std_logic_vector(27 downto 0) := "0000000001110111001100111101";
signal SV14_dim4 : std_logic_vector(27 downto 0) := "0000000000000101101101011100";
signal SV14_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111111101100";
signal SV14_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011000110011";
signal SV14_dim7 : std_logic_vector(27 downto 0) := "0000000000011000111100001010";
signal SV15_dim0 : std_logic_vector(27 downto 0) := "0001000111011101010101010010";
signal SV15_dim1 : std_logic_vector(27 downto 0) := "0000000000000111100000000000";
signal SV15_dim2 : std_logic_vector(27 downto 0) := "0000000010011000011100011111";
signal SV15_dim3 : std_logic_vector(27 downto 0) := "0000000010000011011000010100";
signal SV15_dim4 : std_logic_vector(27 downto 0) := "0000000010100111101100011111";
signal SV15_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101100101001";
signal SV15_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111010111";
signal SV15_dim7 : std_logic_vector(27 downto 0) := "0000000000000101000100101001";
signal SV16_dim0 : std_logic_vector(27 downto 0) := "0000111010111010001101011100";
signal SV16_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101011110110";
signal SV16_dim2 : std_logic_vector(27 downto 0) := "0000000001111010101010101110";
signal SV16_dim3 : std_logic_vector(27 downto 0) := "0000000010001010110000011111";
signal SV16_dim4 : std_logic_vector(27 downto 0) := "0000000000101000110100110011";
signal SV16_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100000000";
signal SV16_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101001001000";
signal SV16_dim7 : std_logic_vector(27 downto 0) := "0000000000001010110110111000";
signal SV17_dim0 : std_logic_vector(27 downto 0) := "0010110011101100000000000000";
signal SV17_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV17_dim2 : std_logic_vector(27 downto 0) := "0000000011100110000000000000";
signal SV17_dim3 : std_logic_vector(27 downto 0) := "0000000010001010000001001000";
signal SV17_dim4 : std_logic_vector(27 downto 0) := "0000000001110100011101001000";
signal SV17_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010011010111";
signal SV17_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111010111";
signal SV17_dim7 : std_logic_vector(27 downto 0) := "0000000000000110011001010010";
signal SV18_dim0 : std_logic_vector(27 downto 0) := "0000110101010011101000010100";
signal SV18_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101011110110";
signal SV18_dim2 : std_logic_vector(27 downto 0) := "0000000001101111000000000000";
signal SV18_dim3 : std_logic_vector(27 downto 0) := "0000000010010011010000011111";
signal SV18_dim4 : std_logic_vector(27 downto 0) := "0000000000101000110100110011";
signal SV18_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100000000";
signal SV18_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101001001000";
signal SV18_dim7 : std_logic_vector(27 downto 0) := "0000000000001011100001011100";
signal SV19_dim0 : std_logic_vector(27 downto 0) := "0010101001100010000000000000";
signal SV19_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV19_dim2 : std_logic_vector(27 downto 0) := "0000000011011001000000000000";
signal SV19_dim3 : std_logic_vector(27 downto 0) := "0000000010000011010001001000";
signal SV19_dim4 : std_logic_vector(27 downto 0) := "0000000001110100011101001000";
signal SV19_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010011010111";
signal SV19_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111010111";
signal SV19_dim7 : std_logic_vector(27 downto 0) := "0000000000000110000101010010";
signal SV20_dim0 : std_logic_vector(27 downto 0) := "0001011010101000000000000000";
signal SV20_dim1 : std_logic_vector(27 downto 0) := "0000000000000101000000000000";
signal SV20_dim2 : std_logic_vector(27 downto 0) := "0000000100100010000000000000";
signal SV20_dim3 : std_logic_vector(27 downto 0) := "0000000010010001100100001010";
signal SV20_dim4 : std_logic_vector(27 downto 0) := "0000000000000011101111001101";
signal SV20_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100000000";
signal SV20_dim6 : std_logic_vector(27 downto 0) := "0000000000000001000011010111";
signal SV20_dim7 : std_logic_vector(27 downto 0) := "0000000000100101101001100110";
signal SV21_dim0 : std_logic_vector(27 downto 0) := "0001011111101000000000000000";
signal SV21_dim1 : std_logic_vector(27 downto 0) := "0000000000000111100000000000";
signal SV21_dim2 : std_logic_vector(27 downto 0) := "0000000011001100000000000000";
signal SV21_dim3 : std_logic_vector(27 downto 0) := "0000000010000111111000010100";
signal SV21_dim4 : std_logic_vector(27 downto 0) := "0000000010100111101100011111";
signal SV21_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101100101001";
signal SV21_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111010111";
signal SV21_dim7 : std_logic_vector(27 downto 0) := "0000000000000101001111110110";
signal SV22_dim0 : std_logic_vector(27 downto 0) := "0001110101001100000000000000";
signal SV22_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV22_dim2 : std_logic_vector(27 downto 0) := "0000000010010110000000000000";
signal SV22_dim3 : std_logic_vector(27 downto 0) := "0000000010001101011011010111";
signal SV22_dim4 : std_logic_vector(27 downto 0) := "0000000001101011001001001000";
signal SV22_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010110001111";
signal SV22_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101111000011";
signal SV22_dim7 : std_logic_vector(27 downto 0) := "0000000000000110110101010010";
signal SV23_dim0 : std_logic_vector(27 downto 0) := "0001000111100111010101010010";
signal SV23_dim1 : std_logic_vector(27 downto 0) := "0000000000000101000000000000";
signal SV23_dim2 : std_logic_vector(27 downto 0) := "0000000011100101001010101110";
signal SV23_dim3 : std_logic_vector(27 downto 0) := "0000000010010010000100010100";
signal SV23_dim4 : std_logic_vector(27 downto 0) := "0000000000000100111100111101";
signal SV23_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000011100001";
signal SV23_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101101111011";
signal SV23_dim7 : std_logic_vector(27 downto 0) := "0000000000100000110100001010";
signal SV24_dim0 : std_logic_vector(27 downto 0) := "0000001011001110111110001111";
signal SV24_dim1 : std_logic_vector(27 downto 0) := "0000000000000011110110101110";
signal SV24_dim2 : std_logic_vector(27 downto 0) := "0000000000101110100111100001";
signal SV24_dim3 : std_logic_vector(27 downto 0) := "0000000001110001110000010100";
signal SV24_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000001011100";
signal SV24_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000001110001";
signal SV24_dim6 : std_logic_vector(27 downto 0) := "0000000000000000110001011100";
signal SV24_dim7 : std_logic_vector(27 downto 0) := "0000000101110011101101010010";
signal SV25_dim0 : std_logic_vector(27 downto 0) := "0000001011011110001000000000";
signal SV25_dim1 : std_logic_vector(27 downto 0) := "0000000000000011111011010111";
signal SV25_dim2 : std_logic_vector(27 downto 0) := "0000000000101110101110111000";
signal SV25_dim3 : std_logic_vector(27 downto 0) := "0000000001110111010001010010";
signal SV25_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000001001000";
signal SV25_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111110000101";
signal SV25_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101000111101";
signal SV25_dim7 : std_logic_vector(27 downto 0) := "0000000110111101010110101110";
signal SV26_dim0 : std_logic_vector(27 downto 0) := "0001010010101011101010000101";
signal SV26_dim1 : std_logic_vector(27 downto 0) := "0000000000001010000110000101";
signal SV26_dim2 : std_logic_vector(27 downto 0) := "0000000010000010101010101110";
signal SV26_dim3 : std_logic_vector(27 downto 0) := "0000000010000111000011101100";
signal SV26_dim4 : std_logic_vector(27 downto 0) := "0000000100100001000101001000";
signal SV26_dim5 : std_logic_vector(27 downto 0) := "0000000000000000001011110110";
signal SV26_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011010101110";
signal SV26_dim7 : std_logic_vector(27 downto 0) := "0000000000000011111110001111";
signal SV27_dim0 : std_logic_vector(27 downto 0) := "0001000010010010111101111011";
signal SV27_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101001100110";
signal SV27_dim2 : std_logic_vector(27 downto 0) := "0000000010001010101010101110";
signal SV27_dim3 : std_logic_vector(27 downto 0) := "0000000010010011110111010111";
signal SV27_dim4 : std_logic_vector(27 downto 0) := "0000000000101110000111100001";
signal SV27_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110000110011";
signal SV27_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110011010";
signal SV27_dim7 : std_logic_vector(27 downto 0) := "0000000000001010111000110011";
signal SV28_dim0 : std_logic_vector(27 downto 0) := "0000000110110101010010011010";
signal SV28_dim1 : std_logic_vector(27 downto 0) := "0000000000000011111111010111";
signal SV28_dim2 : std_logic_vector(27 downto 0) := "0000000000011011011001100110";
signal SV28_dim3 : std_logic_vector(27 downto 0) := "0000000001111010110001111011";
signal SV28_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000000110011";
signal SV28_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110000101";
signal SV28_dim6 : std_logic_vector(27 downto 0) := "0000000000000000110001011100";
signal SV28_dim7 : std_logic_vector(27 downto 0) := "0000001000010101100100000000";
signal SV29_dim0 : std_logic_vector(27 downto 0) := "0000000101101010010101011100";
signal SV29_dim1 : std_logic_vector(27 downto 0) := "0000000000000011111010111000";
signal SV29_dim2 : std_logic_vector(27 downto 0) := "0000000000010111000111010111";
signal SV29_dim3 : std_logic_vector(27 downto 0) := "0000000001110100100000110011";
signal SV29_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000000011111";
signal SV29_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111111000011";
signal SV29_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100110011";
signal SV29_dim7 : std_logic_vector(27 downto 0) := "0000001010110101011110111000";
signal SV30_dim0 : std_logic_vector(27 downto 0) := "0001101001110111001001111011";
signal SV30_dim1 : std_logic_vector(27 downto 0) := "0000000000001000100011100001";
signal SV30_dim2 : std_logic_vector(27 downto 0) := "0000000011000110000000000000";
signal SV30_dim3 : std_logic_vector(27 downto 0) := "0000000001111010110000000000";
signal SV30_dim4 : std_logic_vector(27 downto 0) := "0000000000101011111110101110";
signal SV30_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100011111";
signal SV30_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101010101110";
signal SV30_dim7 : std_logic_vector(27 downto 0) := "0000000000001001010000010100";
signal SV31_dim0 : std_logic_vector(27 downto 0) := "0001010000001111011010101110";
signal SV31_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101001100110";
signal SV31_dim2 : std_logic_vector(27 downto 0) := "0000000010100111110101010010";
signal SV31_dim3 : std_logic_vector(27 downto 0) := "0000000010010000000111110110";
signal SV31_dim4 : std_logic_vector(27 downto 0) := "0000000000110001000110111000";
signal SV31_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110011100001";
signal SV31_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011001110001";
signal SV31_dim7 : std_logic_vector(27 downto 0) := "0000000000001010010010000101";
signal SV32_dim0 : std_logic_vector(27 downto 0) := "0010100101010101100101001000";
signal SV32_dim1 : std_logic_vector(27 downto 0) := "0000000000000111110111110110";
signal SV32_dim2 : std_logic_vector(27 downto 0) := "0000000101010000000000000000";
signal SV32_dim3 : std_logic_vector(27 downto 0) := "0000000001110111100010011010";
signal SV32_dim4 : std_logic_vector(27 downto 0) := "0000000000101011010010011010";
signal SV32_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010100101001";
signal SV32_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101010101110";
signal SV32_dim7 : std_logic_vector(27 downto 0) := "0000000000001001000101011100";
signal SV33_dim0 : std_logic_vector(27 downto 0) := "0001110100100000101010111000";
signal SV33_dim1 : std_logic_vector(27 downto 0) := "0000000000000101000111110110";
signal SV33_dim2 : std_logic_vector(27 downto 0) := "0000000101101100000000000000";
signal SV33_dim3 : std_logic_vector(27 downto 0) := "0000000010010010000100001010";
signal SV33_dim4 : std_logic_vector(27 downto 0) := "0000000000000101000000001010";
signal SV33_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000011001101";
signal SV33_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101110101110";
signal SV33_dim7 : std_logic_vector(27 downto 0) := "0000000000100000101001110001";
signal SV34_dim0 : std_logic_vector(27 downto 0) := "0000111111010110010001110001";
signal SV34_dim1 : std_logic_vector(27 downto 0) := "0000000000000111101001100110";
signal SV34_dim2 : std_logic_vector(27 downto 0) := "0000000010000100100000000000";
signal SV34_dim3 : std_logic_vector(27 downto 0) := "0000000010010110100111010111";
signal SV34_dim4 : std_logic_vector(27 downto 0) := "0000000000101110000111100001";
signal SV34_dim5 : std_logic_vector(27 downto 0) := "1111111111111111110000110011";
signal SV34_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110011010";
signal SV34_dim7 : std_logic_vector(27 downto 0) := "0000000000001011000101110001";
signal SV35_dim0 : std_logic_vector(27 downto 0) := "0001010001111001010010001111";
signal SV35_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101011100001";
signal SV35_dim2 : std_logic_vector(27 downto 0) := "0000000001100111010101010010";
signal SV35_dim3 : std_logic_vector(27 downto 0) := "0000000010000000010100010100";
signal SV35_dim4 : std_logic_vector(27 downto 0) := "0000000111110010001010001111";
signal SV35_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV35_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV35_dim7 : std_logic_vector(27 downto 0) := "0000000000000010111000000000";
signal SV36_dim0 : std_logic_vector(27 downto 0) := "0001111110110011100010011010";
signal SV36_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101011100001";
signal SV36_dim2 : std_logic_vector(27 downto 0) := "0000000010100000000000000000";
signal SV36_dim3 : std_logic_vector(27 downto 0) := "0000000001111000110100010100";
signal SV36_dim4 : std_logic_vector(27 downto 0) := "0000000111110010001010001111";
signal SV36_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV36_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV36_dim7 : std_logic_vector(27 downto 0) := "0000000000000010101101010010";
signal SV37_dim0 : std_logic_vector(27 downto 0) := "0001010111101000101100111101";
signal SV37_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101111110110";
signal SV37_dim2 : std_logic_vector(27 downto 0) := "0000000001101110000000000000";
signal SV37_dim3 : std_logic_vector(27 downto 0) := "0000000010000000010011110110";
signal SV37_dim4 : std_logic_vector(27 downto 0) := "0000000111110000100101001000";
signal SV37_dim5 : std_logic_vector(27 downto 0) := "1111111111111111101111000011";
signal SV37_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV37_dim7 : std_logic_vector(27 downto 0) := "0000000000000010111000010100";
signal SV38_dim0 : std_logic_vector(27 downto 0) := "0001000001010001110001110001";
signal SV38_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100000000000";
signal SV38_dim2 : std_logic_vector(27 downto 0) := "0000000001010011100011100001";
signal SV38_dim3 : std_logic_vector(27 downto 0) := "0000000010001001101011010111";
signal SV38_dim4 : std_logic_vector(27 downto 0) := "0000000001101011001001001000";
signal SV38_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010110001111";
signal SV38_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101111000011";
signal SV38_dim7 : std_logic_vector(27 downto 0) := "0000000000000110101001100110";
signal SV39_dim0 : std_logic_vector(27 downto 0) := "0000001001111010100100000000";
signal SV39_dim1 : std_logic_vector(27 downto 0) := "0000000000000011110000010100";
signal SV39_dim2 : std_logic_vector(27 downto 0) := "0000000000101010001111100001";
signal SV39_dim3 : std_logic_vector(27 downto 0) := "0000000001111011010001011100";
signal SV39_dim4 : std_logic_vector(27 downto 0) := "0000000000000000000000111101";
signal SV39_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111100111101";
signal SV39_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010100100";
signal SV39_dim7 : std_logic_vector(27 downto 0) := "0000000111111100000011100001";
signal SV40_dim0 : std_logic_vector(27 downto 0) := "0010001110111010101010101110";
signal SV40_dim1 : std_logic_vector(27 downto 0) := "0000000000001010000000000000";
signal SV40_dim2 : std_logic_vector(27 downto 0) := "0000000011100100101010101110";
signal SV40_dim3 : std_logic_vector(27 downto 0) := "0000000010001011001011110110";
signal SV40_dim4 : std_logic_vector(27 downto 0) := "0000000100001011111010000101";
signal SV40_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010110111000";
signal SV40_dim6 : std_logic_vector(27 downto 0) := "0000000000000000110000101001";
signal SV40_dim7 : std_logic_vector(27 downto 0) := "0000000000000100010000001010";
signal SV41_dim0 : std_logic_vector(27 downto 0) := "0001101011101110110010100100";
signal SV41_dim1 : std_logic_vector(27 downto 0) := "0000000000000011110010011010";
signal SV41_dim2 : std_logic_vector(27 downto 0) := "0000000111000111001000001010";
signal SV41_dim3 : std_logic_vector(27 downto 0) := "0000000001110100001010101110";
signal SV41_dim4 : std_logic_vector(27 downto 0) := "0000000000000101111010000101";
signal SV41_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000000010100";
signal SV41_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011000000000";
signal SV41_dim7 : std_logic_vector(27 downto 0) := "0000000000010111111001011100";
signal SV42_dim0 : std_logic_vector(27 downto 0) := "0001001111110111000111000011";
signal SV42_dim1 : std_logic_vector(27 downto 0) := "0000000000001010000000000000";
signal SV42_dim2 : std_logic_vector(27 downto 0) := "0000000001111111110001110001";
signal SV42_dim3 : std_logic_vector(27 downto 0) := "0000000010000101011011110110";
signal SV42_dim4 : std_logic_vector(27 downto 0) := "0000000100001011111010000101";
signal SV42_dim5 : std_logic_vector(27 downto 0) := "0000000000000000010110111000";
signal SV42_dim6 : std_logic_vector(27 downto 0) := "0000000000000000110000101001";
signal SV42_dim7 : std_logic_vector(27 downto 0) := "0000000000000100000100110011";
signal SV43_dim0 : std_logic_vector(27 downto 0) := "0001100010011110100111010111";
signal SV43_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101100000000";
signal SV43_dim2 : std_logic_vector(27 downto 0) := "0000000001111100001011110110";
signal SV43_dim3 : std_logic_vector(27 downto 0) := "0000000001111100110010011010";
signal SV43_dim4 : std_logic_vector(27 downto 0) := "0000000000011010001111100001";
signal SV43_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000001110001";
signal SV43_dim6 : std_logic_vector(27 downto 0) := "0000000000000000101100101001";
signal SV43_dim7 : std_logic_vector(27 downto 0) := "0000000000001100001011100001";
signal SV44_dim0 : std_logic_vector(27 downto 0) := "0001101011011011000000000000";
signal SV44_dim1 : std_logic_vector(27 downto 0) := "0000000000001110001100010100";
signal SV44_dim2 : std_logic_vector(27 downto 0) := "0000000001111001000111000011";
signal SV44_dim3 : std_logic_vector(27 downto 0) := "0000000001110110001101110001";
signal SV44_dim4 : std_logic_vector(27 downto 0) := "0000000001010010000110101110";
signal SV44_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000111001101";
signal SV44_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110100100";
signal SV44_dim7 : std_logic_vector(27 downto 0) := "0000000000000110100001011100";
signal SV45_dim0 : std_logic_vector(27 downto 0) := "0001101011100111100000000000";
signal SV45_dim1 : std_logic_vector(27 downto 0) := "0000000000001110011000010100";
signal SV45_dim2 : std_logic_vector(27 downto 0) := "0000000001110111101111100001";
signal SV45_dim3 : std_logic_vector(27 downto 0) := "0000000001101111001110101110";
signal SV45_dim4 : std_logic_vector(27 downto 0) := "0000000000010001101101110001";
signal SV45_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111101100110";
signal SV45_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010011010";
signal SV45_dim7 : std_logic_vector(27 downto 0) := "0000000000001101001101100110";
signal SV46_dim0 : std_logic_vector(27 downto 0) := "0001101010100000111100011111";
signal SV46_dim1 : std_logic_vector(27 downto 0) := "0000000000001111000000111101";
signal SV46_dim2 : std_logic_vector(27 downto 0) := "0000000001110001100000011111";
signal SV46_dim3 : std_logic_vector(27 downto 0) := "0000000001110001001101110001";
signal SV46_dim4 : std_logic_vector(27 downto 0) := "0000000001010010000110101110";
signal SV46_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000111001101";
signal SV46_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110100100";
signal SV46_dim7 : std_logic_vector(27 downto 0) := "0000000000000110001111110110";
signal SV47_dim0 : std_logic_vector(27 downto 0) := "0010111001000000000000000000";
signal SV47_dim1 : std_logic_vector(27 downto 0) := "0000000000001110110001011100";
signal SV47_dim2 : std_logic_vector(27 downto 0) := "0000000011001000011000001010";
signal SV47_dim3 : std_logic_vector(27 downto 0) := "0000000001111111011001010010";
signal SV47_dim4 : std_logic_vector(27 downto 0) := "0000000000011000010111010111";
signal SV47_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110011010";
signal SV47_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100110101110";
signal SV47_dim7 : std_logic_vector(27 downto 0) := "0000000000001100111001111011";
signal SV48_dim0 : std_logic_vector(27 downto 0) := "0001010111010111000111000011";
signal SV48_dim1 : std_logic_vector(27 downto 0) := "0000000000001111000101011100";
signal SV48_dim2 : std_logic_vector(27 downto 0) := "0000000001011100101010001111";
signal SV48_dim3 : std_logic_vector(27 downto 0) := "0000000010001000111001010010";
signal SV48_dim4 : std_logic_vector(27 downto 0) := "0000000000011000010111010111";
signal SV48_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110011010";
signal SV48_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100110101110";
signal SV48_dim7 : std_logic_vector(27 downto 0) := "0000000000001101110111100001";
signal SV49_dim0 : std_logic_vector(27 downto 0) := "0001110111100010000000000000";
signal SV49_dim1 : std_logic_vector(27 downto 0) := "0000000000001110011111001101";
signal SV49_dim2 : std_logic_vector(27 downto 0) := "0000000010000100000000011111";
signal SV49_dim3 : std_logic_vector(27 downto 0) := "0000000010000110000010011010";
signal SV49_dim4 : std_logic_vector(27 downto 0) := "0000000000011000000011000011";
signal SV49_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110001111";
signal SV49_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101001000";
signal SV49_dim7 : std_logic_vector(27 downto 0) := "0000000000001101101010101110";
signal SV50_dim0 : std_logic_vector(27 downto 0) := "0010001101001110010101010010";
signal SV50_dim1 : std_logic_vector(27 downto 0) := "0000000000001111111000101001";
signal SV50_dim2 : std_logic_vector(27 downto 0) := "0000000010001110010000001010";
signal SV50_dim3 : std_logic_vector(27 downto 0) := "0000000001110111100111101100";
signal SV50_dim4 : std_logic_vector(27 downto 0) := "0000000000010001001001111011";
signal SV50_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111100101001";
signal SV50_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010011010";
signal SV50_dim7 : std_logic_vector(27 downto 0) := "0000000000001110011100001010";
signal SV51_dim0 : std_logic_vector(27 downto 0) := "0010001110100000000000000000";
signal SV51_dim1 : std_logic_vector(27 downto 0) := "0000000000001111110111100001";
signal SV51_dim2 : std_logic_vector(27 downto 0) := "0000000010001111101100010100";
signal SV51_dim3 : std_logic_vector(27 downto 0) := "0000000001111101000010011010";
signal SV51_dim4 : std_logic_vector(27 downto 0) := "0000000000011000000011000011";
signal SV51_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110001111";
signal SV51_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101001000";
signal SV51_dim7 : std_logic_vector(27 downto 0) := "0000000000001100110000000000";
signal SV52_dim0 : std_logic_vector(27 downto 0) := "0011000011001011111010001111";
signal SV52_dim1 : std_logic_vector(27 downto 0) := "0000000000001100100001100110";
signal SV52_dim2 : std_logic_vector(27 downto 0) := "0000000011111001010101001000";
signal SV52_dim3 : std_logic_vector(27 downto 0) := "0000000010001110001110100100";
signal SV52_dim4 : std_logic_vector(27 downto 0) := "0000000000011011000110011010";
signal SV52_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110111000";
signal SV52_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100111110110";
signal SV52_dim7 : std_logic_vector(27 downto 0) := "0000000000001101101010001111";
signal SV53_dim0 : std_logic_vector(27 downto 0) := "0001111100101100000000000000";
signal SV53_dim1 : std_logic_vector(27 downto 0) := "0000000000001110010100111101";
signal SV53_dim2 : std_logic_vector(27 downto 0) := "0000000010001011001110111000";
signal SV53_dim3 : std_logic_vector(27 downto 0) := "0000000001111100100100001010";
signal SV53_dim4 : std_logic_vector(27 downto 0) := "0000000000011000010100010100";
signal SV53_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000100010100";
signal SV53_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101001000";
signal SV53_dim7 : std_logic_vector(27 downto 0) := "0000000000001100101000010100";
signal SV54_dim0 : std_logic_vector(27 downto 0) := "0010011001110111001000101001";
signal SV54_dim1 : std_logic_vector(27 downto 0) := "0000000000001011001011101100";
signal SV54_dim2 : std_logic_vector(27 downto 0) := "0000000011011100001000101001";
signal SV54_dim3 : std_logic_vector(27 downto 0) := "0000000001110111111111110110";
signal SV54_dim4 : std_logic_vector(27 downto 0) := "0000000000011000010111010111";
signal SV54_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000111000011";
signal SV54_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101111011";
signal SV54_dim7 : std_logic_vector(27 downto 0) := "0000000000001100001001111011";
signal SV55_dim0 : std_logic_vector(27 downto 0) := "0010111110010100000000000000";
signal SV55_dim1 : std_logic_vector(27 downto 0) := "0000000000001111101001001000";
signal SV55_dim2 : std_logic_vector(27 downto 0) := "0000000011000010101001100110";
signal SV55_dim3 : std_logic_vector(27 downto 0) := "0000000001110111101110101110";
signal SV55_dim4 : std_logic_vector(27 downto 0) := "0000000000010001101101110001";
signal SV55_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111101100110";
signal SV55_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010011010";
signal SV55_dim7 : std_logic_vector(27 downto 0) := "0000000000001110001110001111";
signal SV56_dim0 : std_logic_vector(27 downto 0) := "0001101010010100000000000000";
signal SV56_dim1 : std_logic_vector(27 downto 0) := "0000000000001110011000111101";
signal SV56_dim2 : std_logic_vector(27 downto 0) := "0000000001110110001101010010";
signal SV56_dim3 : std_logic_vector(27 downto 0) := "0000000001111111110100001010";
signal SV56_dim4 : std_logic_vector(27 downto 0) := "0000000000011000010100010100";
signal SV56_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000100010100";
signal SV56_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101001000";
signal SV56_dim7 : std_logic_vector(27 downto 0) := "0000000000001100111101011100";
signal SV57_dim0 : std_logic_vector(27 downto 0) := "0010110010000100000000000000";
signal SV57_dim1 : std_logic_vector(27 downto 0) := "0000000000001111001100010100";
signal SV57_dim2 : std_logic_vector(27 downto 0) := "0000000010111011100000111101";
signal SV57_dim3 : std_logic_vector(27 downto 0) := "0000000010000110011110111000";
signal SV57_dim4 : std_logic_vector(27 downto 0) := "0000000000011001011100111101";
signal SV57_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110111000";
signal SV57_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100111101";
signal SV57_dim7 : std_logic_vector(27 downto 0) := "0000000000001101010100111101";
signal SV58_dim0 : std_logic_vector(27 downto 0) := "0001010001100110100000001010";
signal SV58_dim1 : std_logic_vector(27 downto 0) := "0000000000001011010110000101";
signal SV58_dim2 : std_logic_vector(27 downto 0) := "0000000001110011000101001000";
signal SV58_dim3 : std_logic_vector(27 downto 0) := "0000000001101010010110011010";
signal SV58_dim4 : std_logic_vector(27 downto 0) := "0000000000010011010100010100";
signal SV58_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111110011010";
signal SV58_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100001110001";
signal SV58_dim7 : std_logic_vector(27 downto 0) := "0000000000001100000110011010";
signal SV59_dim0 : std_logic_vector(27 downto 0) := "0001001100110101110110100100";
signal SV59_dim1 : std_logic_vector(27 downto 0) := "0000000000001011011110101110";
signal SV59_dim2 : std_logic_vector(27 downto 0) := "0000000001101011000110001111";
signal SV59_dim3 : std_logic_vector(27 downto 0) := "0000000001101101100110111000";
signal SV59_dim4 : std_logic_vector(27 downto 0) := "0000000000011010001111001101";
signal SV59_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111111110110";
signal SV59_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100000000";
signal SV59_dim7 : std_logic_vector(27 downto 0) := "0000000000001010101100110011";
signal SV60_dim0 : std_logic_vector(27 downto 0) := "0001110010101110100000000000";
signal SV60_dim1 : std_logic_vector(27 downto 0) := "0000000000001111010110101110";
signal SV60_dim2 : std_logic_vector(27 downto 0) := "0000000001110111100010011010";
signal SV60_dim3 : std_logic_vector(27 downto 0) := "0000000001111011001101110001";
signal SV60_dim4 : std_logic_vector(27 downto 0) := "0000000001010010000110101110";
signal SV60_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000111001101";
signal SV60_dim6 : std_logic_vector(27 downto 0) := "0000000000000000011110100100";
signal SV60_dim7 : std_logic_vector(27 downto 0) := "0000000000000110110011001101";
signal SV61_dim0 : std_logic_vector(27 downto 0) := "0010001011001000101010101110";
signal SV61_dim1 : std_logic_vector(27 downto 0) := "0000000000001101111000000000";
signal SV61_dim2 : std_logic_vector(27 downto 0) := "0000000010100000011101010010";
signal SV61_dim3 : std_logic_vector(27 downto 0) := "0000000010001001001110111000";
signal SV61_dim4 : std_logic_vector(27 downto 0) := "0000000000011001011100111101";
signal SV61_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110111000";
signal SV61_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100111101";
signal SV61_dim7 : std_logic_vector(27 downto 0) := "0000000000001101100110011010";
signal SV62_dim0 : std_logic_vector(27 downto 0) := "0001000001101111101110001111";
signal SV62_dim1 : std_logic_vector(27 downto 0) := "0000000000001110011000011111";
signal SV62_dim2 : std_logic_vector(27 downto 0) := "0000000001001001001001010010";
signal SV62_dim3 : std_logic_vector(27 downto 0) := "0000000001111010010011101100";
signal SV62_dim4 : std_logic_vector(27 downto 0) := "0000000000011000011111010111";
signal SV62_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000100001010";
signal SV62_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100011110110";
signal SV62_dim7 : std_logic_vector(27 downto 0) := "0000000000001100010110111000";
signal SV63_dim0 : std_logic_vector(27 downto 0) := "0001001011001010100001111011";
signal SV63_dim1 : std_logic_vector(27 downto 0) := "0000000000001101001110101110";
signal SV63_dim2 : std_logic_vector(27 downto 0) := "0000000001011010111001110001";
signal SV63_dim3 : std_logic_vector(27 downto 0) := "0000000010000011100100110011";
signal SV63_dim4 : std_logic_vector(27 downto 0) := "0000000000010000101100101001";
signal SV63_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111101011100";
signal SV63_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010111000";
signal SV63_dim7 : std_logic_vector(27 downto 0) := "0000000000010000000110011010";
signal SV64_dim0 : std_logic_vector(27 downto 0) := "0001010110010101010101010010";
signal SV64_dim1 : std_logic_vector(27 downto 0) := "0000000000010000000010000101";
signal SV64_dim2 : std_logic_vector(27 downto 0) := "0000000001010110001001111011";
signal SV64_dim3 : std_logic_vector(27 downto 0) := "0000000010000011101110111000";
signal SV64_dim4 : std_logic_vector(27 downto 0) := "0000000000011001011100111101";
signal SV64_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000110111000";
signal SV64_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100111101";
signal SV64_dim7 : std_logic_vector(27 downto 0) := "0000000000001101000011100001";
signal SV65_dim0 : std_logic_vector(27 downto 0) := "0001011000001010000000000000";
signal SV65_dim1 : std_logic_vector(27 downto 0) := "0000000000001110000111110110";
signal SV65_dim2 : std_logic_vector(27 downto 0) := "0000000001100011110111101100";
signal SV65_dim3 : std_logic_vector(27 downto 0) := "0000000001110000001100111101";
signal SV65_dim4 : std_logic_vector(27 downto 0) := "0000000000011000111000111101";
signal SV65_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000000000000";
signal SV65_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101100110";
signal SV65_dim7 : std_logic_vector(27 downto 0) := "0000000000001011001111101100";
signal SV66_dim0 : std_logic_vector(27 downto 0) := "0001001001000011101010101110";
signal SV66_dim1 : std_logic_vector(27 downto 0) := "0000000000001111011100101001";
signal SV66_dim2 : std_logic_vector(27 downto 0) := "0000000001001011101010101110";
signal SV66_dim3 : std_logic_vector(27 downto 0) := "0000000001110111101100111101";
signal SV66_dim4 : std_logic_vector(27 downto 0) := "0000000000011000111000111101";
signal SV66_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000000000000";
signal SV66_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100101100110";
signal SV66_dim7 : std_logic_vector(27 downto 0) := "0000000000001011111111110110";
signal SV67_dim0 : std_logic_vector(27 downto 0) := "0010101000110101100010101110";
signal SV67_dim1 : std_logic_vector(27 downto 0) := "0000000000001100101100010100";
signal SV67_dim2 : std_logic_vector(27 downto 0) := "0000000011010100110110101110";
signal SV67_dim3 : std_logic_vector(27 downto 0) := "0000000010000100110010111000";
signal SV67_dim4 : std_logic_vector(27 downto 0) := "0000000000011001011001100110";
signal SV67_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000100000000";
signal SV67_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100100101001";
signal SV67_dim7 : std_logic_vector(27 downto 0) := "0000000000001101001011001101";
signal SV68_dim0 : std_logic_vector(27 downto 0) := "0010010100000011010111110110";
signal SV68_dim1 : std_logic_vector(27 downto 0) := "0000000000001011111011101100";
signal SV68_dim2 : std_logic_vector(27 downto 0) := "0000000011000110100000110011";
signal SV68_dim3 : std_logic_vector(27 downto 0) := "0000000010000010010100011111";
signal SV68_dim4 : std_logic_vector(27 downto 0) := "0000000000010111101100010100";
signal SV68_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000011101100";
signal SV68_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100011010111";
signal SV68_dim7 : std_logic_vector(27 downto 0) := "0000000000001101011000110011";
signal SV69_dim0 : std_logic_vector(27 downto 0) := "0010011010010111000000000000";
signal SV69_dim1 : std_logic_vector(27 downto 0) := "0000000000001111011011000011";
signal SV69_dim2 : std_logic_vector(27 downto 0) := "0000000010100000001000101001";
signal SV69_dim3 : std_logic_vector(27 downto 0) := "0000000001110111010011101100";
signal SV69_dim4 : std_logic_vector(27 downto 0) := "0000000000011000011111010111";
signal SV69_dim5 : std_logic_vector(27 downto 0) := "0000000000000000000100001010";
signal SV69_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100011110110";
signal SV69_dim7 : std_logic_vector(27 downto 0) := "0000000000001100000011100001";
signal SV70_dim0 : std_logic_vector(27 downto 0) := "0001100011000101010101010010";
signal SV70_dim1 : std_logic_vector(27 downto 0) := "0000000000001110010111010111";
signal SV70_dim2 : std_logic_vector(27 downto 0) := "0000000001101110010110101110";
signal SV70_dim3 : std_logic_vector(27 downto 0) := "0000000001111110100111101100";
signal SV70_dim4 : std_logic_vector(27 downto 0) := "0000000000010001001001111011";
signal SV70_dim5 : std_logic_vector(27 downto 0) := "1111111111111111111100101001";
signal SV70_dim6 : std_logic_vector(27 downto 0) := "0000000000000000100010011010";
signal SV70_dim7 : std_logic_vector(27 downto 0) := "0000000000001111010010001111";

signal SV0_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV1_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV2_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV3_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV4_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV5_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV6_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV7_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV8_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV9_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV10_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV11_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV12_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV13_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV14_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV15_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV16_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV17_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV18_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV19_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV20_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV21_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV22_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV23_alphaY : std_logic_vector(11 downto 0) := "110101100110";
signal SV24_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV25_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV26_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV27_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV28_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV29_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV30_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV31_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV32_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV33_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV34_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV35_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV36_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV37_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV38_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV39_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV40_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV41_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV42_alphaY : std_logic_vector(11 downto 0) := "110101100101";
signal SV43_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV44_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV45_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV46_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV47_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV48_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV49_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV50_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV51_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV52_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV53_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV54_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV55_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV56_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV57_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV58_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV59_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV60_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV61_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV62_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV63_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV64_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV65_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV66_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV67_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV68_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV69_alphaY : std_logic_vector(11 downto 0) := "010000000000";
signal SV70_alphaY : std_logic_vector(11 downto 0) := "010000000000";

signal gamma : std_logic_vector(11 downto 0) := "010110001110"; --  1.388 1.011000111000111001

signal b : std_logic_vector(19 downto 0) := "11111111111010011011";  -- (-)0.34883721 0.0101100101001101011 ca2(00000000000101100101) 11111111111010011010 + 1 

signal output : std_logic;

signal test_data_dim0 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim1 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim2 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim3 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim4 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim5 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim6 : std_logic_vector(27 downto 0) := (others => '0'); 
signal test_data_dim7 : std_logic_vector(27 downto 0) := (others => '0'); 

begin

	TOP_0 : TOP
		port map(	SV0_dim0 => SV0_dim0,
					SV0_dim1 => SV0_dim1,
					SV0_dim2 => SV0_dim2,
					SV0_dim3 => SV0_dim3,
					SV0_dim4 => SV0_dim4,
					SV0_dim5 => SV0_dim5,
					SV0_dim6 => SV0_dim6,
					SV0_dim7 => SV0_dim7,
					SV1_dim0 => SV1_dim0,
					SV1_dim1 => SV1_dim1,
					SV1_dim2 => SV1_dim2,
					SV1_dim3 => SV1_dim3,
					SV1_dim4 => SV1_dim4,
					SV1_dim5 => SV1_dim5,
					SV1_dim6 => SV1_dim6,
					SV1_dim7 => SV1_dim7,
					SV2_dim0 => SV2_dim0,
					SV2_dim1 => SV2_dim1,
					SV2_dim2 => SV2_dim2,
					SV2_dim3 => SV2_dim3,
					SV2_dim4 => SV2_dim4,
					SV2_dim5 => SV2_dim5,
					SV2_dim6 => SV2_dim6,
					SV2_dim7 => SV2_dim7,
					SV3_dim0 => SV3_dim0,
					SV3_dim1 => SV3_dim1,
					SV3_dim2 => SV3_dim2,
					SV3_dim3 => SV3_dim3,
					SV3_dim4 => SV3_dim4,
					SV3_dim5 => SV3_dim5,
					SV3_dim6 => SV3_dim6,
					SV3_dim7 => SV3_dim7,
					SV4_dim0 => SV4_dim0,
					SV4_dim1 => SV4_dim1,
					SV4_dim2 => SV4_dim2,
					SV4_dim3 => SV4_dim3,
					SV4_dim4 => SV4_dim4,
					SV4_dim5 => SV4_dim5,
					SV4_dim6 => SV4_dim6,
					SV4_dim7 => SV4_dim7,
					SV5_dim0 => SV5_dim0,
					SV5_dim1 => SV5_dim1,
					SV5_dim2 => SV5_dim2,
					SV5_dim3 => SV5_dim3,
					SV5_dim4 => SV5_dim4,
					SV5_dim5 => SV5_dim5,
					SV5_dim6 => SV5_dim6,
					SV5_dim7 => SV5_dim7,
					SV6_dim0 => SV6_dim0,
					SV6_dim1 => SV6_dim1,
					SV6_dim2 => SV6_dim2,
					SV6_dim3 => SV6_dim3,
					SV6_dim4 => SV6_dim4,
					SV6_dim5 => SV6_dim5,
					SV6_dim6 => SV6_dim6,
					SV6_dim7 => SV6_dim7,
					SV7_dim0 => SV7_dim0,
					SV7_dim1 => SV7_dim1,
					SV7_dim2 => SV7_dim2,
					SV7_dim3 => SV7_dim3,
					SV7_dim4 => SV7_dim4,
					SV7_dim5 => SV7_dim5,
					SV7_dim6 => SV7_dim6,
					SV7_dim7 => SV7_dim7,
					SV8_dim0 => SV8_dim0,
					SV8_dim1 => SV8_dim1,
					SV8_dim2 => SV8_dim2,
					SV8_dim3 => SV8_dim3,
					SV8_dim4 => SV8_dim4,
					SV8_dim5 => SV8_dim5,
					SV8_dim6 => SV8_dim6,
					SV8_dim7 => SV8_dim7,
					SV9_dim0 => SV9_dim0,
					SV9_dim1 => SV9_dim1,
					SV9_dim2 => SV9_dim2,
					SV9_dim3 => SV9_dim3,
					SV9_dim4 => SV9_dim4,
					SV9_dim5 => SV9_dim5,
					SV9_dim6 => SV9_dim6,
					SV9_dim7 => SV9_dim7,
					SV10_dim0 => SV10_dim0,
					SV10_dim1 => SV10_dim1,
					SV10_dim2 => SV10_dim2,
					SV10_dim3 => SV10_dim3,
					SV10_dim4 => SV10_dim4,
					SV10_dim5 => SV10_dim5,
					SV10_dim6 => SV10_dim6,
					SV10_dim7 => SV10_dim7,
					SV11_dim0 => SV11_dim0,
					SV11_dim1 => SV11_dim1,
					SV11_dim2 => SV11_dim2,
					SV11_dim3 => SV11_dim3,
					SV11_dim4 => SV11_dim4,
					SV11_dim5 => SV11_dim5,
					SV11_dim6 => SV11_dim6,
					SV11_dim7 => SV11_dim7,
					SV12_dim0 => SV12_dim0,
					SV12_dim1 => SV12_dim1,
					SV12_dim2 => SV12_dim2,
					SV12_dim3 => SV12_dim3,
					SV12_dim4 => SV12_dim4,
					SV12_dim5 => SV12_dim5,
					SV12_dim6 => SV12_dim6,
					SV12_dim7 => SV12_dim7,
					SV13_dim0 => SV13_dim0,
					SV13_dim1 => SV13_dim1,
					SV13_dim2 => SV13_dim2,
					SV13_dim3 => SV13_dim3,
					SV13_dim4 => SV13_dim4,
					SV13_dim5 => SV13_dim5,
					SV13_dim6 => SV13_dim6,
					SV13_dim7 => SV13_dim7,
					SV14_dim0 => SV14_dim0,
					SV14_dim1 => SV14_dim1,
					SV14_dim2 => SV14_dim2,
					SV14_dim3 => SV14_dim3,
					SV14_dim4 => SV14_dim4,
					SV14_dim5 => SV14_dim5,
					SV14_dim6 => SV14_dim6,
					SV14_dim7 => SV14_dim7,
					SV15_dim0 => SV15_dim0,
					SV15_dim1 => SV15_dim1,
					SV15_dim2 => SV15_dim2,
					SV15_dim3 => SV15_dim3,
					SV15_dim4 => SV15_dim4,
					SV15_dim5 => SV15_dim5,
					SV15_dim6 => SV15_dim6,
					SV15_dim7 => SV15_dim7,
					SV16_dim0 => SV16_dim0,
					SV16_dim1 => SV16_dim1,
					SV16_dim2 => SV16_dim2,
					SV16_dim3 => SV16_dim3,
					SV16_dim4 => SV16_dim4,
					SV16_dim5 => SV16_dim5,
					SV16_dim6 => SV16_dim6,
					SV16_dim7 => SV16_dim7,
					SV17_dim0 => SV17_dim0,
					SV17_dim1 => SV17_dim1,
					SV17_dim2 => SV17_dim2,
					SV17_dim3 => SV17_dim3,
					SV17_dim4 => SV17_dim4,
					SV17_dim5 => SV17_dim5,
					SV17_dim6 => SV17_dim6,
					SV17_dim7 => SV17_dim7,
					SV18_dim0 => SV18_dim0,
					SV18_dim1 => SV18_dim1,
					SV18_dim2 => SV18_dim2,
					SV18_dim3 => SV18_dim3,
					SV18_dim4 => SV18_dim4,
					SV18_dim5 => SV18_dim5,
					SV18_dim6 => SV18_dim6,
					SV18_dim7 => SV18_dim7,
					SV19_dim0 => SV19_dim0,
					SV19_dim1 => SV19_dim1,
					SV19_dim2 => SV19_dim2,
					SV19_dim3 => SV19_dim3,
					SV19_dim4 => SV19_dim4,
					SV19_dim5 => SV19_dim5,
					SV19_dim6 => SV19_dim6,
					SV19_dim7 => SV19_dim7,
					SV20_dim0 => SV20_dim0,
					SV20_dim1 => SV20_dim1,
					SV20_dim2 => SV20_dim2,
					SV20_dim3 => SV20_dim3,
					SV20_dim4 => SV20_dim4,
					SV20_dim5 => SV20_dim5,
					SV20_dim6 => SV20_dim6,
					SV20_dim7 => SV20_dim7,
					SV21_dim0 => SV21_dim0,
					SV21_dim1 => SV21_dim1,
					SV21_dim2 => SV21_dim2,
					SV21_dim3 => SV21_dim3,
					SV21_dim4 => SV21_dim4,
					SV21_dim5 => SV21_dim5,
					SV21_dim6 => SV21_dim6,
					SV21_dim7 => SV21_dim7,
					SV22_dim0 => SV22_dim0,
					SV22_dim1 => SV22_dim1,
					SV22_dim2 => SV22_dim2,
					SV22_dim3 => SV22_dim3,
					SV22_dim4 => SV22_dim4,
					SV22_dim5 => SV22_dim5,
					SV22_dim6 => SV22_dim6,
					SV22_dim7 => SV22_dim7,
					SV23_dim0 => SV23_dim0,
					SV23_dim1 => SV23_dim1,
					SV23_dim2 => SV23_dim2,
					SV23_dim3 => SV23_dim3,
					SV23_dim4 => SV23_dim4,
					SV23_dim5 => SV23_dim5,
					SV23_dim6 => SV23_dim6,
					SV23_dim7 => SV23_dim7,
					SV24_dim0 => SV24_dim0,
					SV24_dim1 => SV24_dim1,
					SV24_dim2 => SV24_dim2,
					SV24_dim3 => SV24_dim3,
					SV24_dim4 => SV24_dim4,
					SV24_dim5 => SV24_dim5,
					SV24_dim6 => SV24_dim6,
					SV24_dim7 => SV24_dim7,
					SV25_dim0 => SV25_dim0,
					SV25_dim1 => SV25_dim1,
					SV25_dim2 => SV25_dim2,
					SV25_dim3 => SV25_dim3,
					SV25_dim4 => SV25_dim4,
					SV25_dim5 => SV25_dim5,
					SV25_dim6 => SV25_dim6,
					SV25_dim7 => SV25_dim7,
					SV26_dim0 => SV26_dim0,
					SV26_dim1 => SV26_dim1,
					SV26_dim2 => SV26_dim2,
					SV26_dim3 => SV26_dim3,
					SV26_dim4 => SV26_dim4,
					SV26_dim5 => SV26_dim5,
					SV26_dim6 => SV26_dim6,
					SV26_dim7 => SV26_dim7,
					SV27_dim0 => SV27_dim0,
					SV27_dim1 => SV27_dim1,
					SV27_dim2 => SV27_dim2,
					SV27_dim3 => SV27_dim3,
					SV27_dim4 => SV27_dim4,
					SV27_dim5 => SV27_dim5,
					SV27_dim6 => SV27_dim6,
					SV27_dim7 => SV27_dim7,
					SV28_dim0 => SV28_dim0,
					SV28_dim1 => SV28_dim1,
					SV28_dim2 => SV28_dim2,
					SV28_dim3 => SV28_dim3,
					SV28_dim4 => SV28_dim4,
					SV28_dim5 => SV28_dim5,
					SV28_dim6 => SV28_dim6,
					SV28_dim7 => SV28_dim7,
					SV29_dim0 => SV29_dim0,
					SV29_dim1 => SV29_dim1,
					SV29_dim2 => SV29_dim2,
					SV29_dim3 => SV29_dim3,
					SV29_dim4 => SV29_dim4,
					SV29_dim5 => SV29_dim5,
					SV29_dim6 => SV29_dim6,
					SV29_dim7 => SV29_dim7,
					SV30_dim0 => SV30_dim0,
					SV30_dim1 => SV30_dim1,
					SV30_dim2 => SV30_dim2,
					SV30_dim3 => SV30_dim3,
					SV30_dim4 => SV30_dim4,
					SV30_dim5 => SV30_dim5,
					SV30_dim6 => SV30_dim6,
					SV30_dim7 => SV30_dim7,
					SV31_dim0 => SV31_dim0,
					SV31_dim1 => SV31_dim1,
					SV31_dim2 => SV31_dim2,
					SV31_dim3 => SV31_dim3,
					SV31_dim4 => SV31_dim4,
					SV31_dim5 => SV31_dim5,
					SV31_dim6 => SV31_dim6,
					SV31_dim7 => SV31_dim7,
					SV32_dim0 => SV32_dim0,
					SV32_dim1 => SV32_dim1,
					SV32_dim2 => SV32_dim2,
					SV32_dim3 => SV32_dim3,
					SV32_dim4 => SV32_dim4,
					SV32_dim5 => SV32_dim5,
					SV32_dim6 => SV32_dim6,
					SV32_dim7 => SV32_dim7,
					SV33_dim0 => SV33_dim0,
					SV33_dim1 => SV33_dim1,
					SV33_dim2 => SV33_dim2,
					SV33_dim3 => SV33_dim3,
					SV33_dim4 => SV33_dim4,
					SV33_dim5 => SV33_dim5,
					SV33_dim6 => SV33_dim6,
					SV33_dim7 => SV33_dim7,
					SV34_dim0 => SV34_dim0,
					SV34_dim1 => SV34_dim1,
					SV34_dim2 => SV34_dim2,
					SV34_dim3 => SV34_dim3,
					SV34_dim4 => SV34_dim4,
					SV34_dim5 => SV34_dim5,
					SV34_dim6 => SV34_dim6,
					SV34_dim7 => SV34_dim7,
					SV35_dim0 => SV35_dim0,
					SV35_dim1 => SV35_dim1,
					SV35_dim2 => SV35_dim2,
					SV35_dim3 => SV35_dim3,
					SV35_dim4 => SV35_dim4,
					SV35_dim5 => SV35_dim5,
					SV35_dim6 => SV35_dim6,
					SV35_dim7 => SV35_dim7,
					SV36_dim0 => SV36_dim0,
					SV36_dim1 => SV36_dim1,
					SV36_dim2 => SV36_dim2,
					SV36_dim3 => SV36_dim3,
					SV36_dim4 => SV36_dim4,
					SV36_dim5 => SV36_dim5,
					SV36_dim6 => SV36_dim6,
					SV36_dim7 => SV36_dim7,
					SV37_dim0 => SV37_dim0,
					SV37_dim1 => SV37_dim1,
					SV37_dim2 => SV37_dim2,
					SV37_dim3 => SV37_dim3,
					SV37_dim4 => SV37_dim4,
					SV37_dim5 => SV37_dim5,
					SV37_dim6 => SV37_dim6,
					SV37_dim7 => SV37_dim7,
					SV38_dim0 => SV38_dim0,
					SV38_dim1 => SV38_dim1,
					SV38_dim2 => SV38_dim2,
					SV38_dim3 => SV38_dim3,
					SV38_dim4 => SV38_dim4,
					SV38_dim5 => SV38_dim5,
					SV38_dim6 => SV38_dim6,
					SV38_dim7 => SV38_dim7,
					SV39_dim0 => SV39_dim0,
					SV39_dim1 => SV39_dim1,
					SV39_dim2 => SV39_dim2,
					SV39_dim3 => SV39_dim3,
					SV39_dim4 => SV39_dim4,
					SV39_dim5 => SV39_dim5,
					SV39_dim6 => SV39_dim6,
					SV39_dim7 => SV39_dim7,
					SV40_dim0 => SV40_dim0,
					SV40_dim1 => SV40_dim1,
					SV40_dim2 => SV40_dim2,
					SV40_dim3 => SV40_dim3,
					SV40_dim4 => SV40_dim4,
					SV40_dim5 => SV40_dim5,
					SV40_dim6 => SV40_dim6,
					SV40_dim7 => SV40_dim7,
					SV41_dim0 => SV41_dim0,
					SV41_dim1 => SV41_dim1,
					SV41_dim2 => SV41_dim2,
					SV41_dim3 => SV41_dim3,
					SV41_dim4 => SV41_dim4,
					SV41_dim5 => SV41_dim5,
					SV41_dim6 => SV41_dim6,
					SV41_dim7 => SV41_dim7,
					SV42_dim0 => SV42_dim0,
					SV42_dim1 => SV42_dim1,
					SV42_dim2 => SV42_dim2,
					SV42_dim3 => SV42_dim3,
					SV42_dim4 => SV42_dim4,
					SV42_dim5 => SV42_dim5,
					SV42_dim6 => SV42_dim6,
					SV42_dim7 => SV42_dim7,
					SV43_dim0 => SV43_dim0,
					SV43_dim1 => SV43_dim1,
					SV43_dim2 => SV43_dim2,
					SV43_dim3 => SV43_dim3,
					SV43_dim4 => SV43_dim4,
					SV43_dim5 => SV43_dim5,
					SV43_dim6 => SV43_dim6,
					SV43_dim7 => SV43_dim7,
					SV44_dim0 => SV44_dim0,
					SV44_dim1 => SV44_dim1,
					SV44_dim2 => SV44_dim2,
					SV44_dim3 => SV44_dim3,
					SV44_dim4 => SV44_dim4,
					SV44_dim5 => SV44_dim5,
					SV44_dim6 => SV44_dim6,
					SV44_dim7 => SV44_dim7,
					SV45_dim0 => SV45_dim0,
					SV45_dim1 => SV45_dim1,
					SV45_dim2 => SV45_dim2,
					SV45_dim3 => SV45_dim3,
					SV45_dim4 => SV45_dim4,
					SV45_dim5 => SV45_dim5,
					SV45_dim6 => SV45_dim6,
					SV45_dim7 => SV45_dim7,
					SV46_dim0 => SV46_dim0,
					SV46_dim1 => SV46_dim1,
					SV46_dim2 => SV46_dim2,
					SV46_dim3 => SV46_dim3,
					SV46_dim4 => SV46_dim4,
					SV46_dim5 => SV46_dim5,
					SV46_dim6 => SV46_dim6,
					SV46_dim7 => SV46_dim7,
					SV47_dim0 => SV47_dim0,
					SV47_dim1 => SV47_dim1,
					SV47_dim2 => SV47_dim2,
					SV47_dim3 => SV47_dim3,
					SV47_dim4 => SV47_dim4,
					SV47_dim5 => SV47_dim5,
					SV47_dim6 => SV47_dim6,
					SV47_dim7 => SV47_dim7,
					SV48_dim0 => SV48_dim0,
					SV48_dim1 => SV48_dim1,
					SV48_dim2 => SV48_dim2,
					SV48_dim3 => SV48_dim3,
					SV48_dim4 => SV48_dim4,
					SV48_dim5 => SV48_dim5,
					SV48_dim6 => SV48_dim6,
					SV48_dim7 => SV48_dim7,
					SV49_dim0 => SV49_dim0,
					SV49_dim1 => SV49_dim1,
					SV49_dim2 => SV49_dim2,
					SV49_dim3 => SV49_dim3,
					SV49_dim4 => SV49_dim4,
					SV49_dim5 => SV49_dim5,
					SV49_dim6 => SV49_dim6,
					SV49_dim7 => SV49_dim7,
					SV50_dim0 => SV50_dim0,
					SV50_dim1 => SV50_dim1,
					SV50_dim2 => SV50_dim2,
					SV50_dim3 => SV50_dim3,
					SV50_dim4 => SV50_dim4,
					SV50_dim5 => SV50_dim5,
					SV50_dim6 => SV50_dim6,
					SV50_dim7 => SV50_dim7,
					SV51_dim0 => SV51_dim0,
					SV51_dim1 => SV51_dim1,
					SV51_dim2 => SV51_dim2,
					SV51_dim3 => SV51_dim3,
					SV51_dim4 => SV51_dim4,
					SV51_dim5 => SV51_dim5,
					SV51_dim6 => SV51_dim6,
					SV51_dim7 => SV51_dim7,
					SV52_dim0 => SV52_dim0,
					SV52_dim1 => SV52_dim1,
					SV52_dim2 => SV52_dim2,
					SV52_dim3 => SV52_dim3,
					SV52_dim4 => SV52_dim4,
					SV52_dim5 => SV52_dim5,
					SV52_dim6 => SV52_dim6,
					SV52_dim7 => SV52_dim7,
					SV53_dim0 => SV53_dim0,
					SV53_dim1 => SV53_dim1,
					SV53_dim2 => SV53_dim2,
					SV53_dim3 => SV53_dim3,
					SV53_dim4 => SV53_dim4,
					SV53_dim5 => SV53_dim5,
					SV53_dim6 => SV53_dim6,
					SV53_dim7 => SV53_dim7,
					SV54_dim0 => SV54_dim0,
					SV54_dim1 => SV54_dim1,
					SV54_dim2 => SV54_dim2,
					SV54_dim3 => SV54_dim3,
					SV54_dim4 => SV54_dim4,
					SV54_dim5 => SV54_dim5,
					SV54_dim6 => SV54_dim6,
					SV54_dim7 => SV54_dim7,
					SV55_dim0 => SV55_dim0,
					SV55_dim1 => SV55_dim1,
					SV55_dim2 => SV55_dim2,
					SV55_dim3 => SV55_dim3,
					SV55_dim4 => SV55_dim4,
					SV55_dim5 => SV55_dim5,
					SV55_dim6 => SV55_dim6,
					SV55_dim7 => SV55_dim7,
					SV56_dim0 => SV56_dim0,
					SV56_dim1 => SV56_dim1,
					SV56_dim2 => SV56_dim2,
					SV56_dim3 => SV56_dim3,
					SV56_dim4 => SV56_dim4,
					SV56_dim5 => SV56_dim5,
					SV56_dim6 => SV56_dim6,
					SV56_dim7 => SV56_dim7,
					SV57_dim0 => SV57_dim0,
					SV57_dim1 => SV57_dim1,
					SV57_dim2 => SV57_dim2,
					SV57_dim3 => SV57_dim3,
					SV57_dim4 => SV57_dim4,
					SV57_dim5 => SV57_dim5,
					SV57_dim6 => SV57_dim6,
					SV57_dim7 => SV57_dim7,
					SV58_dim0 => SV58_dim0,
					SV58_dim1 => SV58_dim1,
					SV58_dim2 => SV58_dim2,
					SV58_dim3 => SV58_dim3,
					SV58_dim4 => SV58_dim4,
					SV58_dim5 => SV58_dim5,
					SV58_dim6 => SV58_dim6,
					SV58_dim7 => SV58_dim7,
					SV59_dim0 => SV59_dim0,
					SV59_dim1 => SV59_dim1,
					SV59_dim2 => SV59_dim2,
					SV59_dim3 => SV59_dim3,
					SV59_dim4 => SV59_dim4,
					SV59_dim5 => SV59_dim5,
					SV59_dim6 => SV59_dim6,
					SV59_dim7 => SV59_dim7,
					SV60_dim0 => SV60_dim0,
					SV60_dim1 => SV60_dim1,
					SV60_dim2 => SV60_dim2,
					SV60_dim3 => SV60_dim3,
					SV60_dim4 => SV60_dim4,
					SV60_dim5 => SV60_dim5,
					SV60_dim6 => SV60_dim6,
					SV60_dim7 => SV60_dim7,
					SV61_dim0 => SV61_dim0,
					SV61_dim1 => SV61_dim1,
					SV61_dim2 => SV61_dim2,
					SV61_dim3 => SV61_dim3,
					SV61_dim4 => SV61_dim4,
					SV61_dim5 => SV61_dim5,
					SV61_dim6 => SV61_dim6,
					SV61_dim7 => SV61_dim7,
					SV62_dim0 => SV62_dim0,
					SV62_dim1 => SV62_dim1,
					SV62_dim2 => SV62_dim2,
					SV62_dim3 => SV62_dim3,
					SV62_dim4 => SV62_dim4,
					SV62_dim5 => SV62_dim5,
					SV62_dim6 => SV62_dim6,
					SV62_dim7 => SV62_dim7,
					SV63_dim0 => SV63_dim0,
					SV63_dim1 => SV63_dim1,
					SV63_dim2 => SV63_dim2,
					SV63_dim3 => SV63_dim3,
					SV63_dim4 => SV63_dim4,
					SV63_dim5 => SV63_dim5,
					SV63_dim6 => SV63_dim6,
					SV63_dim7 => SV63_dim7,
					SV64_dim0 => SV64_dim0,
					SV64_dim1 => SV64_dim1,
					SV64_dim2 => SV64_dim2,
					SV64_dim3 => SV64_dim3,
					SV64_dim4 => SV64_dim4,
					SV64_dim5 => SV64_dim5,
					SV64_dim6 => SV64_dim6,
					SV64_dim7 => SV64_dim7,
					SV65_dim0 => SV65_dim0,
					SV65_dim1 => SV65_dim1,
					SV65_dim2 => SV65_dim2,
					SV65_dim3 => SV65_dim3,
					SV65_dim4 => SV65_dim4,
					SV65_dim5 => SV65_dim5,
					SV65_dim6 => SV65_dim6,
					SV65_dim7 => SV65_dim7,
					SV66_dim0 => SV66_dim0,
					SV66_dim1 => SV66_dim1,
					SV66_dim2 => SV66_dim2,
					SV66_dim3 => SV66_dim3,
					SV66_dim4 => SV66_dim4,
					SV66_dim5 => SV66_dim5,
					SV66_dim6 => SV66_dim6,
					SV66_dim7 => SV66_dim7,
					SV67_dim0 => SV67_dim0,
					SV67_dim1 => SV67_dim1,
					SV67_dim2 => SV67_dim2,
					SV67_dim3 => SV67_dim3,
					SV67_dim4 => SV67_dim4,
					SV67_dim5 => SV67_dim5,
					SV67_dim6 => SV67_dim6,
					SV67_dim7 => SV67_dim7,
					SV68_dim0 => SV68_dim0,
					SV68_dim1 => SV68_dim1,
					SV68_dim2 => SV68_dim2,
					SV68_dim3 => SV68_dim3,
					SV68_dim4 => SV68_dim4,
					SV68_dim5 => SV68_dim5,
					SV68_dim6 => SV68_dim6,
					SV68_dim7 => SV68_dim7,
					SV69_dim0 => SV69_dim0,
					SV69_dim1 => SV69_dim1,
					SV69_dim2 => SV69_dim2,
					SV69_dim3 => SV69_dim3,
					SV69_dim4 => SV69_dim4,
					SV69_dim5 => SV69_dim5,
					SV69_dim6 => SV69_dim6,
					SV69_dim7 => SV69_dim7,
					SV70_dim0 => SV70_dim0,
					SV70_dim1 => SV70_dim1,
					SV70_dim2 => SV70_dim2,
					SV70_dim3 => SV70_dim3,
					SV70_dim4 => SV70_dim4,
					SV70_dim5 => SV70_dim5,
					SV70_dim6 => SV70_dim6,
					SV70_dim7 => SV70_dim7,
					test_data_dim0 => test_data_dim0, 
					test_data_dim1 => test_data_dim1, 
					test_data_dim2 => test_data_dim2, 
					test_data_dim3 => test_data_dim3, 
					test_data_dim4 => test_data_dim4, 
					test_data_dim5 => test_data_dim5, 
					test_data_dim6 => test_data_dim6, 
					test_data_dim7 => test_data_dim7, 
					SV0_alphaY => SV0_alphaY, 
					SV1_alphaY => SV1_alphaY, 
					SV2_alphaY => SV2_alphaY, 
					SV3_alphaY => SV3_alphaY, 
					SV4_alphaY => SV4_alphaY, 
					SV5_alphaY => SV5_alphaY, 
					SV6_alphaY => SV6_alphaY, 
					SV7_alphaY => SV7_alphaY, 
					SV8_alphaY => SV8_alphaY, 
					SV9_alphaY => SV9_alphaY, 
					SV10_alphaY => SV10_alphaY, 
					SV11_alphaY => SV11_alphaY, 
					SV12_alphaY => SV12_alphaY, 
					SV13_alphaY => SV13_alphaY, 
					SV14_alphaY => SV14_alphaY, 
					SV15_alphaY => SV15_alphaY, 
					SV16_alphaY => SV16_alphaY, 
					SV17_alphaY => SV17_alphaY, 
					SV18_alphaY => SV18_alphaY, 
					SV19_alphaY => SV19_alphaY, 
					SV20_alphaY => SV20_alphaY, 
					SV21_alphaY => SV21_alphaY, 
					SV22_alphaY => SV22_alphaY, 
					SV23_alphaY => SV23_alphaY, 
					SV24_alphaY => SV24_alphaY, 
					SV25_alphaY => SV25_alphaY, 
					SV26_alphaY => SV26_alphaY, 
					SV27_alphaY => SV27_alphaY, 
					SV28_alphaY => SV28_alphaY, 
					SV29_alphaY => SV29_alphaY, 
					SV30_alphaY => SV30_alphaY, 
					SV31_alphaY => SV31_alphaY, 
					SV32_alphaY => SV32_alphaY, 
					SV33_alphaY => SV33_alphaY, 
					SV34_alphaY => SV34_alphaY, 
					SV35_alphaY => SV35_alphaY, 
					SV36_alphaY => SV36_alphaY, 
					SV37_alphaY => SV37_alphaY, 
					SV38_alphaY => SV38_alphaY, 
					SV39_alphaY => SV39_alphaY, 
					SV40_alphaY => SV40_alphaY, 
					SV41_alphaY => SV41_alphaY, 
					SV42_alphaY => SV42_alphaY, 
					SV43_alphaY => SV43_alphaY, 
					SV44_alphaY => SV44_alphaY, 
					SV45_alphaY => SV45_alphaY, 
					SV46_alphaY => SV46_alphaY, 
					SV47_alphaY => SV47_alphaY, 
					SV48_alphaY => SV48_alphaY, 
					SV49_alphaY => SV49_alphaY, 
					SV50_alphaY => SV50_alphaY, 
					SV51_alphaY => SV51_alphaY, 
					SV52_alphaY => SV52_alphaY, 
					SV53_alphaY => SV53_alphaY, 
					SV54_alphaY => SV54_alphaY, 
					SV55_alphaY => SV55_alphaY, 
					SV56_alphaY => SV56_alphaY, 
					SV57_alphaY => SV57_alphaY, 
					SV58_alphaY => SV58_alphaY, 
					SV59_alphaY => SV59_alphaY, 
					SV60_alphaY => SV60_alphaY, 
					SV61_alphaY => SV61_alphaY, 
					SV62_alphaY => SV62_alphaY, 
					SV63_alphaY => SV63_alphaY, 
					SV64_alphaY => SV64_alphaY, 
					SV65_alphaY => SV65_alphaY, 
					SV66_alphaY => SV66_alphaY, 
					SV67_alphaY => SV67_alphaY, 
					SV68_alphaY => SV68_alphaY, 
					SV69_alphaY => SV69_alphaY, 
					SV70_alphaY => SV70_alphaY, 
					gamma => gamma, 
					b => b, 
					output => output 
					);
					
	test_data_dim0 <= "0001101101110111111101110001" after 10 ns, "0010100100000001100000000000" after 20 ns, "0000110111111100000000010100" after 30 ns, "0001010100101001100110101110" after 40 ns, "0010011101110101000000000000" after 50 ns, "0001011101011100101101111011" after 60 ns, "0001011001010101110101010010" after 70 ns, "0010111001101000000000000000" after 80 ns, "0010000011000110110001001000" after 90 ns, "0001101000010100100101100110" after 100 ns, "0001111000011010101010101110" after 110 ns, "0001010011001100000110111000" after 120 ns, "0001001011001011001011101100" after 130 ns, "0000111111010011100110011010" after 140 ns, "0000001000100011100110000101" after 150 ns, "0010101111111101101000001010" after 160 ns, "0000111110001010100110101110" after 170 ns, "0010100111010110000000000000" after 180 ns;
	test_data_dim1 <= "0000000000000100100101011100" after 10 ns, "0000000000001111010111101100" after 20 ns, "0000000000000111101001100110" after 30 ns, "0000000000001100100110011010" after 40 ns, "0000000000010000001101011100" after 50 ns, "0000000000001100101111100001" after 60 ns, "0000000000001111001000001010" after 70 ns, "0000000000000111100000000000" after 80 ns, "0000000000000111101011110110" after 90 ns, "0000000000001010000110000101" after 100 ns, "0000000000001010000000000000" after 110 ns, "0000000000000111101001100110" after 120 ns, "0000000000001000100101111011" after 130 ns, "0000000000000100110000010100" after 140 ns, "0000000000000011110000000000" after 150 ns, "0000000000001010001111001101" after 160 ns, "0000000000000100100111101100" after 170 ns, "0000000000001110111000000000" after 180 ns;
	test_data_dim2 <= "0000000101111111100000000000" after 10 ns, "0000000010101010101111000011" after 20 ns, "0000000001110101000000000000" after 30 ns, "0000000001101011100000000000" after 40 ns, "0000000010011011110001110001" after 50 ns, "0000000001110101010101010010" after 60 ns, "0000000001011110011111100001" after 70 ns, "0000000110001100000000000000" after 80 ns, "0000000100010001000000000000" after 90 ns, "0000000010100101010101010010" after 100 ns, "0000000011000000101010101110" after 110 ns, "0000000010101110000000000000" after 120 ns, "0000000010001100000000000000" after 130 ns, "0000000011010101000000000000" after 140 ns, "0000000000100100011111110110" after 150 ns, "0000000100010011000000000000" after 160 ns, "0000000011010111010101010010" after 170 ns, "0000000010110100000000010100" after 180 ns;
	test_data_dim3 <= "0000000001110101010110101110" after 10 ns, "0000000001111010100000011111" after 20 ns, "0000000010010110100111110110" after 30 ns, "0000000001111100101010011010" after 40 ns, "0000000001111101010100001010" after 50 ns, "0000000010000001111010101110" after 60 ns, "0000000001110010100000011111" after 70 ns, "0000000001111100011000010100" after 80 ns, "0000000010010000010000011111" after 90 ns, "0000000010001101000011101100" after 100 ns, "0000000010001110011011110110" after 110 ns, "0000000010010011101000010100" after 120 ns, "0000000001110101110000000000" after 130 ns, "0000000001101111010101110001" after 140 ns, "0000000001100111101111001101" after 150 ns, "0000000010000011010001010010" after 160 ns, "0000000001110010010101111011" after 170 ns, "0000000001111001010100001010" after 180 ns;
	test_data_dim4 <= "0000000000000111100010100100" after 10 ns, "0000000000011001000011110110" after 20 ns, "0000000000110001000110111000" after 30 ns, "0000000010010111101110000101" after 40 ns, "0000000000011000011111010111" after 50 ns, "0000000010010111010011010111" after 60 ns, "0000000000011001000011110110" after 70 ns, "0000000010100111101100011111" after 80 ns, "0000000000101000110100110011" after 90 ns, "0000000100100001000101001000" after 100 ns, "0000000100001011111010000101" after 110 ns, "0000000000110000110100101001" after 120 ns, "0000000000101100000000010100" after 130 ns, "0000000000000111101110101110" after 140 ns, "0000000000000000000001011100" after 150 ns, "0000000001011111011110111000" after 160 ns, "0000000000000111101010101110" after 170 ns, "0000000000011000010100010100" after 180 ns;
	test_data_dim5 <= "1111111111111111111101110001" after 10 ns, "0000000000000000000001100110" after 20 ns, "1111111111111111110011100001" after 30 ns, "0000000000000000000111000011" after 40 ns, "0000000000000000000100001010" after 50 ns, "0000000000000000000111000011" after 60 ns, "0000000000000000000001100110" after 70 ns, "1111111111111111101100101001" after 80 ns, "0000000000000000010100000000" after 90 ns, "0000000000000000001011110110" after 100 ns, "0000000000000000010110111000" after 110 ns, "1111111111111111110011010111" after 120 ns, "0000000000000000010100011111" after 130 ns, "1111111111111111111101110001" after 140 ns, "0000000000000000000000010100" after 150 ns, "0000000000000000001000000000" after 160 ns, "1111111111111111111101110001" after 170 ns, "0000000000000000000100010100" after 180 ns;
	test_data_dim6 <= "0000000000000000011111110110" after 10 ns, "0000000000000000100100111101" after 20 ns, "0000000000000000011001110001" after 30 ns, "0000000000000000010011000011" after 40 ns, "0000000000000000100011110110" after 50 ns, "0000000000000000010011000011" after 60 ns, "0000000000000000100100111101" after 70 ns, "0000000000000000100111010111" after 80 ns, "0000000000000000101001001000" after 90 ns, "0000000000000000011010101110" after 100 ns, "0000000000000000110000101001" after 110 ns, "0000000000000000011001111011" after 120 ns, "0000000000000000101010101110" after 130 ns, "0000000000000000100000010100" after 140 ns, "0000000000000000101011001101" after 150 ns, "0000000000000000010100000000" after 160 ns, "0000000000000000100000000000" after 170 ns, "0000000000000000100101001000" after 180 ns;
	test_data_dim7 <= "0000000000010101010111101100" after 10 ns, "0000000000001100001111000011" after 20 ns, "0000000000001010101111110110" after 30 ns, "0000000000000101000011110110" after 40 ns, "0000000000001100101010001111" after 50 ns, "0000000000000101010001111011" after 60 ns, "0000000000001011011100000000" after 70 ns, "0000000000000100110011010111" after 80 ns, "0000000000001011010010011010" after 90 ns, "0000000000000100001001011100" after 100 ns, "0000000000000100010110011010" after 110 ns, "0000000000001010100100001010" after 120 ns, "0000000000001000111000000000" after 130 ns, "0000000000010100000001011100" after 140 ns, "0000000101010100110000000000" after 150 ns, "0000000000000110101101111011" after 160 ns, "0000000000010100101001011100" after 170 ns, "0000000000001100010011001101" after 180 ns;


end Behavioral;
