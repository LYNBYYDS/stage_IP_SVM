Mon Drive
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 
-- Design Name: 
-- Module Name: TOP - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TOP is
    Port (  -- SV
            SV0_dim0 : in std_logic_vector(27 downto 0); 
            SV0_dim1 : in std_logic_vector(27 downto 0); 
            SV0_dim2 : in std_logic_vector(27 downto 0); 
            SV0_dim3 : in std_logic_vector(27 downto 0); 
            SV0_dim4 : in std_logic_vector(27 downto 0); 
            SV0_dim5 : in std_logic_vector(27 downto 0); 
            SV0_dim6 : in std_logic_vector(27 downto 0); 
            SV0_dim7 : in std_logic_vector(27 downto 0); 
            SV1_dim0 : in std_logic_vector(27 downto 0); 
            SV1_dim1 : in std_logic_vector(27 downto 0); 
            SV1_dim2 : in std_logic_vector(27 downto 0); 
            SV1_dim3 : in std_logic_vector(27 downto 0); 
            SV1_dim4 : in std_logic_vector(27 downto 0); 
            SV1_dim5 : in std_logic_vector(27 downto 0); 
            SV1_dim6 : in std_logic_vector(27 downto 0); 
            SV1_dim7 : in std_logic_vector(27 downto 0); 
            SV2_dim0 : in std_logic_vector(27 downto 0); 
            SV2_dim1 : in std_logic_vector(27 downto 0); 
            SV2_dim2 : in std_logic_vector(27 downto 0); 
            SV2_dim3 : in std_logic_vector(27 downto 0); 
            SV2_dim4 : in std_logic_vector(27 downto 0); 
            SV2_dim5 : in std_logic_vector(27 downto 0); 
            SV2_dim6 : in std_logic_vector(27 downto 0); 
            SV2_dim7 : in std_logic_vector(27 downto 0); 
            SV3_dim0 : in std_logic_vector(27 downto 0); 
            SV3_dim1 : in std_logic_vector(27 downto 0); 
            SV3_dim2 : in std_logic_vector(27 downto 0); 
            SV3_dim3 : in std_logic_vector(27 downto 0); 
            SV3_dim4 : in std_logic_vector(27 downto 0); 
            SV3_dim5 : in std_logic_vector(27 downto 0); 
            SV3_dim6 : in std_logic_vector(27 downto 0); 
            SV3_dim7 : in std_logic_vector(27 downto 0); 
            SV4_dim0 : in std_logic_vector(27 downto 0); 
            SV4_dim1 : in std_logic_vector(27 downto 0); 
            SV4_dim2 : in std_logic_vector(27 downto 0); 
            SV4_dim3 : in std_logic_vector(27 downto 0); 
            SV4_dim4 : in std_logic_vector(27 downto 0); 
            SV4_dim5 : in std_logic_vector(27 downto 0); 
            SV4_dim6 : in std_logic_vector(27 downto 0); 
            SV4_dim7 : in std_logic_vector(27 downto 0); 
            SV5_dim0 : in std_logic_vector(27 downto 0); 
            SV5_dim1 : in std_logic_vector(27 downto 0); 
            SV5_dim2 : in std_logic_vector(27 downto 0); 
            SV5_dim3 : in std_logic_vector(27 downto 0); 
            SV5_dim4 : in std_logic_vector(27 downto 0); 
            SV5_dim5 : in std_logic_vector(27 downto 0); 
            SV5_dim6 : in std_logic_vector(27 downto 0); 
            SV5_dim7 : in std_logic_vector(27 downto 0); 
            SV6_dim0 : in std_logic_vector(27 downto 0); 
            SV6_dim1 : in std_logic_vector(27 downto 0); 
            SV6_dim2 : in std_logic_vector(27 downto 0); 
            SV6_dim3 : in std_logic_vector(27 downto 0); 
            SV6_dim4 : in std_logic_vector(27 downto 0); 
            SV6_dim5 : in std_logic_vector(27 downto 0); 
            SV6_dim6 : in std_logic_vector(27 downto 0); 
            SV6_dim7 : in std_logic_vector(27 downto 0); 
            SV7_dim0 : in std_logic_vector(27 downto 0); 
            SV7_dim1 : in std_logic_vector(27 downto 0); 
            SV7_dim2 : in std_logic_vector(27 downto 0); 
            SV7_dim3 : in std_logic_vector(27 downto 0); 
            SV7_dim4 : in std_logic_vector(27 downto 0); 
            SV7_dim5 : in std_logic_vector(27 downto 0); 
            SV7_dim6 : in std_logic_vector(27 downto 0); 
            SV7_dim7 : in std_logic_vector(27 downto 0); 
            SV8_dim0 : in std_logic_vector(27 downto 0); 
            SV8_dim1 : in std_logic_vector(27 downto 0); 
            SV8_dim2 : in std_logic_vector(27 downto 0); 
            SV8_dim3 : in std_logic_vector(27 downto 0); 
            SV8_dim4 : in std_logic_vector(27 downto 0); 
            SV8_dim5 : in std_logic_vector(27 downto 0); 
            SV8_dim6 : in std_logic_vector(27 downto 0); 
            SV8_dim7 : in std_logic_vector(27 downto 0); 
            SV9_dim0 : in std_logic_vector(27 downto 0); 
            SV9_dim1 : in std_logic_vector(27 downto 0); 
            SV9_dim2 : in std_logic_vector(27 downto 0); 
            SV9_dim3 : in std_logic_vector(27 downto 0); 
            SV9_dim4 : in std_logic_vector(27 downto 0); 
            SV9_dim5 : in std_logic_vector(27 downto 0); 
            SV9_dim6 : in std_logic_vector(27 downto 0); 
            SV9_dim7 : in std_logic_vector(27 downto 0); 
            SV10_dim0 : in std_logic_vector(27 downto 0); 
            SV10_dim1 : in std_logic_vector(27 downto 0); 
            SV10_dim2 : in std_logic_vector(27 downto 0); 
            SV10_dim3 : in std_logic_vector(27 downto 0); 
            SV10_dim4 : in std_logic_vector(27 downto 0); 
            SV10_dim5 : in std_logic_vector(27 downto 0); 
            SV10_dim6 : in std_logic_vector(27 downto 0); 
            SV10_dim7 : in std_logic_vector(27 downto 0); 
            SV11_dim0 : in std_logic_vector(27 downto 0); 
            SV11_dim1 : in std_logic_vector(27 downto 0); 
            SV11_dim2 : in std_logic_vector(27 downto 0); 
            SV11_dim3 : in std_logic_vector(27 downto 0); 
            SV11_dim4 : in std_logic_vector(27 downto 0); 
            SV11_dim5 : in std_logic_vector(27 downto 0); 
            SV11_dim6 : in std_logic_vector(27 downto 0); 
            SV11_dim7 : in std_logic_vector(27 downto 0); 
            SV12_dim0 : in std_logic_vector(27 downto 0); 
            SV12_dim1 : in std_logic_vector(27 downto 0); 
            SV12_dim2 : in std_logic_vector(27 downto 0); 
            SV12_dim3 : in std_logic_vector(27 downto 0); 
            SV12_dim4 : in std_logic_vector(27 downto 0); 
            SV12_dim5 : in std_logic_vector(27 downto 0); 
            SV12_dim6 : in std_logic_vector(27 downto 0); 
            SV12_dim7 : in std_logic_vector(27 downto 0); 
            SV13_dim0 : in std_logic_vector(27 downto 0); 
            SV13_dim1 : in std_logic_vector(27 downto 0); 
            SV13_dim2 : in std_logic_vector(27 downto 0); 
            SV13_dim3 : in std_logic_vector(27 downto 0); 
            SV13_dim4 : in std_logic_vector(27 downto 0); 
            SV13_dim5 : in std_logic_vector(27 downto 0); 
            SV13_dim6 : in std_logic_vector(27 downto 0); 
            SV13_dim7 : in std_logic_vector(27 downto 0); 
            SV14_dim0 : in std_logic_vector(27 downto 0); 
            SV14_dim1 : in std_logic_vector(27 downto 0); 
            SV14_dim2 : in std_logic_vector(27 downto 0); 
            SV14_dim3 : in std_logic_vector(27 downto 0); 
            SV14_dim4 : in std_logic_vector(27 downto 0); 
            SV14_dim5 : in std_logic_vector(27 downto 0); 
            SV14_dim6 : in std_logic_vector(27 downto 0); 
            SV14_dim7 : in std_logic_vector(27 downto 0); 
            SV15_dim0 : in std_logic_vector(27 downto 0); 
            SV15_dim1 : in std_logic_vector(27 downto 0); 
            SV15_dim2 : in std_logic_vector(27 downto 0); 
            SV15_dim3 : in std_logic_vector(27 downto 0); 
            SV15_dim4 : in std_logic_vector(27 downto 0); 
            SV15_dim5 : in std_logic_vector(27 downto 0); 
            SV15_dim6 : in std_logic_vector(27 downto 0); 
            SV15_dim7 : in std_logic_vector(27 downto 0); 
            SV16_dim0 : in std_logic_vector(27 downto 0); 
            SV16_dim1 : in std_logic_vector(27 downto 0); 
            SV16_dim2 : in std_logic_vector(27 downto 0); 
            SV16_dim3 : in std_logic_vector(27 downto 0); 
            SV16_dim4 : in std_logic_vector(27 downto 0); 
            SV16_dim5 : in std_logic_vector(27 downto 0); 
            SV16_dim6 : in std_logic_vector(27 downto 0); 
            SV16_dim7 : in std_logic_vector(27 downto 0); 
            SV17_dim0 : in std_logic_vector(27 downto 0); 
            SV17_dim1 : in std_logic_vector(27 downto 0); 
            SV17_dim2 : in std_logic_vector(27 downto 0); 
            SV17_dim3 : in std_logic_vector(27 downto 0); 
            SV17_dim4 : in std_logic_vector(27 downto 0); 
            SV17_dim5 : in std_logic_vector(27 downto 0); 
            SV17_dim6 : in std_logic_vector(27 downto 0); 
            SV17_dim7 : in std_logic_vector(27 downto 0); 
            SV18_dim0 : in std_logic_vector(27 downto 0); 
            SV18_dim1 : in std_logic_vector(27 downto 0); 
            SV18_dim2 : in std_logic_vector(27 downto 0); 
            SV18_dim3 : in std_logic_vector(27 downto 0); 
            SV18_dim4 : in std_logic_vector(27 downto 0); 
            SV18_dim5 : in std_logic_vector(27 downto 0); 
            SV18_dim6 : in std_logic_vector(27 downto 0); 
            SV18_dim7 : in std_logic_vector(27 downto 0); 
            SV19_dim0 : in std_logic_vector(27 downto 0); 
            SV19_dim1 : in std_logic_vector(27 downto 0); 
            SV19_dim2 : in std_logic_vector(27 downto 0); 
            SV19_dim3 : in std_logic_vector(27 downto 0); 
            SV19_dim4 : in std_logic_vector(27 downto 0); 
            SV19_dim5 : in std_logic_vector(27 downto 0); 
            SV19_dim6 : in std_logic_vector(27 downto 0); 
            SV19_dim7 : in std_logic_vector(27 downto 0); 
            SV20_dim0 : in std_logic_vector(27 downto 0); 
            SV20_dim1 : in std_logic_vector(27 downto 0); 
            SV20_dim2 : in std_logic_vector(27 downto 0); 
            SV20_dim3 : in std_logic_vector(27 downto 0); 
            SV20_dim4 : in std_logic_vector(27 downto 0); 
            SV20_dim5 : in std_logic_vector(27 downto 0); 
            SV20_dim6 : in std_logic_vector(27 downto 0); 
            SV20_dim7 : in std_logic_vector(27 downto 0); 
            SV21_dim0 : in std_logic_vector(27 downto 0); 
            SV21_dim1 : in std_logic_vector(27 downto 0); 
            SV21_dim2 : in std_logic_vector(27 downto 0); 
            SV21_dim3 : in std_logic_vector(27 downto 0); 
            SV21_dim4 : in std_logic_vector(27 downto 0); 
            SV21_dim5 : in std_logic_vector(27 downto 0); 
            SV21_dim6 : in std_logic_vector(27 downto 0); 
            SV21_dim7 : in std_logic_vector(27 downto 0); 
            SV22_dim0 : in std_logic_vector(27 downto 0); 
            SV22_dim1 : in std_logic_vector(27 downto 0); 
            SV22_dim2 : in std_logic_vector(27 downto 0); 
            SV22_dim3 : in std_logic_vector(27 downto 0); 
            SV22_dim4 : in std_logic_vector(27 downto 0); 
            SV22_dim5 : in std_logic_vector(27 downto 0); 
            SV22_dim6 : in std_logic_vector(27 downto 0); 
            SV22_dim7 : in std_logic_vector(27 downto 0); 
            SV23_dim0 : in std_logic_vector(27 downto 0); 
            SV23_dim1 : in std_logic_vector(27 downto 0); 
            SV23_dim2 : in std_logic_vector(27 downto 0); 
            SV23_dim3 : in std_logic_vector(27 downto 0); 
            SV23_dim4 : in std_logic_vector(27 downto 0); 
            SV23_dim5 : in std_logic_vector(27 downto 0); 
            SV23_dim6 : in std_logic_vector(27 downto 0); 
            SV23_dim7 : in std_logic_vector(27 downto 0); 
            SV24_dim0 : in std_logic_vector(27 downto 0); 
            SV24_dim1 : in std_logic_vector(27 downto 0); 
            SV24_dim2 : in std_logic_vector(27 downto 0); 
            SV24_dim3 : in std_logic_vector(27 downto 0); 
            SV24_dim4 : in std_logic_vector(27 downto 0); 
            SV24_dim5 : in std_logic_vector(27 downto 0); 
            SV24_dim6 : in std_logic_vector(27 downto 0); 
            SV24_dim7 : in std_logic_vector(27 downto 0); 
            SV25_dim0 : in std_logic_vector(27 downto 0); 
            SV25_dim1 : in std_logic_vector(27 downto 0); 
            SV25_dim2 : in std_logic_vector(27 downto 0); 
            SV25_dim3 : in std_logic_vector(27 downto 0); 
            SV25_dim4 : in std_logic_vector(27 downto 0); 
            SV25_dim5 : in std_logic_vector(27 downto 0); 
            SV25_dim6 : in std_logic_vector(27 downto 0); 
            SV25_dim7 : in std_logic_vector(27 downto 0); 
            SV26_dim0 : in std_logic_vector(27 downto 0); 
            SV26_dim1 : in std_logic_vector(27 downto 0); 
            SV26_dim2 : in std_logic_vector(27 downto 0); 
            SV26_dim3 : in std_logic_vector(27 downto 0); 
            SV26_dim4 : in std_logic_vector(27 downto 0); 
            SV26_dim5 : in std_logic_vector(27 downto 0); 
            SV26_dim6 : in std_logic_vector(27 downto 0); 
            SV26_dim7 : in std_logic_vector(27 downto 0); 
            SV27_dim0 : in std_logic_vector(27 downto 0); 
            SV27_dim1 : in std_logic_vector(27 downto 0); 
            SV27_dim2 : in std_logic_vector(27 downto 0); 
            SV27_dim3 : in std_logic_vector(27 downto 0); 
            SV27_dim4 : in std_logic_vector(27 downto 0); 
            SV27_dim5 : in std_logic_vector(27 downto 0); 
            SV27_dim6 : in std_logic_vector(27 downto 0); 
            SV27_dim7 : in std_logic_vector(27 downto 0); 
            SV28_dim0 : in std_logic_vector(27 downto 0); 
            SV28_dim1 : in std_logic_vector(27 downto 0); 
            SV28_dim2 : in std_logic_vector(27 downto 0); 
            SV28_dim3 : in std_logic_vector(27 downto 0); 
            SV28_dim4 : in std_logic_vector(27 downto 0); 
            SV28_dim5 : in std_logic_vector(27 downto 0); 
            SV28_dim6 : in std_logic_vector(27 downto 0); 
            SV28_dim7 : in std_logic_vector(27 downto 0); 
            SV29_dim0 : in std_logic_vector(27 downto 0); 
            SV29_dim1 : in std_logic_vector(27 downto 0); 
            SV29_dim2 : in std_logic_vector(27 downto 0); 
            SV29_dim3 : in std_logic_vector(27 downto 0); 
            SV29_dim4 : in std_logic_vector(27 downto 0); 
            SV29_dim5 : in std_logic_vector(27 downto 0); 
            SV29_dim6 : in std_logic_vector(27 downto 0); 
            SV29_dim7 : in std_logic_vector(27 downto 0); 
            SV30_dim0 : in std_logic_vector(27 downto 0); 
            SV30_dim1 : in std_logic_vector(27 downto 0); 
            SV30_dim2 : in std_logic_vector(27 downto 0); 
            SV30_dim3 : in std_logic_vector(27 downto 0); 
            SV30_dim4 : in std_logic_vector(27 downto 0); 
            SV30_dim5 : in std_logic_vector(27 downto 0); 
            SV30_dim6 : in std_logic_vector(27 downto 0); 
            SV30_dim7 : in std_logic_vector(27 downto 0); 
            SV31_dim0 : in std_logic_vector(27 downto 0); 
            SV31_dim1 : in std_logic_vector(27 downto 0); 
            SV31_dim2 : in std_logic_vector(27 downto 0); 
            SV31_dim3 : in std_logic_vector(27 downto 0); 
            SV31_dim4 : in std_logic_vector(27 downto 0); 
            SV31_dim5 : in std_logic_vector(27 downto 0); 
            SV31_dim6 : in std_logic_vector(27 downto 0); 
            SV31_dim7 : in std_logic_vector(27 downto 0); 
            SV32_dim0 : in std_logic_vector(27 downto 0); 
            SV32_dim1 : in std_logic_vector(27 downto 0); 
            SV32_dim2 : in std_logic_vector(27 downto 0); 
            SV32_dim3 : in std_logic_vector(27 downto 0); 
            SV32_dim4 : in std_logic_vector(27 downto 0); 
            SV32_dim5 : in std_logic_vector(27 downto 0); 
            SV32_dim6 : in std_logic_vector(27 downto 0); 
            SV32_dim7 : in std_logic_vector(27 downto 0); 
            SV33_dim0 : in std_logic_vector(27 downto 0); 
            SV33_dim1 : in std_logic_vector(27 downto 0); 
            SV33_dim2 : in std_logic_vector(27 downto 0); 
            SV33_dim3 : in std_logic_vector(27 downto 0); 
            SV33_dim4 : in std_logic_vector(27 downto 0); 
            SV33_dim5 : in std_logic_vector(27 downto 0); 
            SV33_dim6 : in std_logic_vector(27 downto 0); 
            SV33_dim7 : in std_logic_vector(27 downto 0); 
            SV34_dim0 : in std_logic_vector(27 downto 0); 
            SV34_dim1 : in std_logic_vector(27 downto 0); 
            SV34_dim2 : in std_logic_vector(27 downto 0); 
            SV34_dim3 : in std_logic_vector(27 downto 0); 
            SV34_dim4 : in std_logic_vector(27 downto 0); 
            SV34_dim5 : in std_logic_vector(27 downto 0); 
            SV34_dim6 : in std_logic_vector(27 downto 0); 
            SV34_dim7 : in std_logic_vector(27 downto 0); 
            SV35_dim0 : in std_logic_vector(27 downto 0); 
            SV35_dim1 : in std_logic_vector(27 downto 0); 
            SV35_dim2 : in std_logic_vector(27 downto 0); 
            SV35_dim3 : in std_logic_vector(27 downto 0); 
            SV35_dim4 : in std_logic_vector(27 downto 0); 
            SV35_dim5 : in std_logic_vector(27 downto 0); 
            SV35_dim6 : in std_logic_vector(27 downto 0); 
            SV35_dim7 : in std_logic_vector(27 downto 0); 
            SV36_dim0 : in std_logic_vector(27 downto 0); 
            SV36_dim1 : in std_logic_vector(27 downto 0); 
            SV36_dim2 : in std_logic_vector(27 downto 0); 
            SV36_dim3 : in std_logic_vector(27 downto 0); 
            SV36_dim4 : in std_logic_vector(27 downto 0); 
            SV36_dim5 : in std_logic_vector(27 downto 0); 
            SV36_dim6 : in std_logic_vector(27 downto 0); 
            SV36_dim7 : in std_logic_vector(27 downto 0); 
            SV37_dim0 : in std_logic_vector(27 downto 0); 
            SV37_dim1 : in std_logic_vector(27 downto 0); 
            SV37_dim2 : in std_logic_vector(27 downto 0); 
            SV37_dim3 : in std_logic_vector(27 downto 0); 
            SV37_dim4 : in std_logic_vector(27 downto 0); 
            SV37_dim5 : in std_logic_vector(27 downto 0); 
            SV37_dim6 : in std_logic_vector(27 downto 0); 
            SV37_dim7 : in std_logic_vector(27 downto 0); 
            SV38_dim0 : in std_logic_vector(27 downto 0); 
            SV38_dim1 : in std_logic_vector(27 downto 0); 
            SV38_dim2 : in std_logic_vector(27 downto 0); 
            SV38_dim3 : in std_logic_vector(27 downto 0); 
            SV38_dim4 : in std_logic_vector(27 downto 0); 
            SV38_dim5 : in std_logic_vector(27 downto 0); 
            SV38_dim6 : in std_logic_vector(27 downto 0); 
            SV38_dim7 : in std_logic_vector(27 downto 0); 
            SV39_dim0 : in std_logic_vector(27 downto 0); 
            SV39_dim1 : in std_logic_vector(27 downto 0); 
            SV39_dim2 : in std_logic_vector(27 downto 0); 
            SV39_dim3 : in std_logic_vector(27 downto 0); 
            SV39_dim4 : in std_logic_vector(27 downto 0); 
            SV39_dim5 : in std_logic_vector(27 downto 0); 
            SV39_dim6 : in std_logic_vector(27 downto 0); 
            SV39_dim7 : in std_logic_vector(27 downto 0); 
            SV40_dim0 : in std_logic_vector(27 downto 0); 
            SV40_dim1 : in std_logic_vector(27 downto 0); 
            SV40_dim2 : in std_logic_vector(27 downto 0); 
            SV40_dim3 : in std_logic_vector(27 downto 0); 
            SV40_dim4 : in std_logic_vector(27 downto 0); 
            SV40_dim5 : in std_logic_vector(27 downto 0); 
            SV40_dim6 : in std_logic_vector(27 downto 0); 
            SV40_dim7 : in std_logic_vector(27 downto 0); 
            SV41_dim0 : in std_logic_vector(27 downto 0); 
            SV41_dim1 : in std_logic_vector(27 downto 0); 
            SV41_dim2 : in std_logic_vector(27 downto 0); 
            SV41_dim3 : in std_logic_vector(27 downto 0); 
            SV41_dim4 : in std_logic_vector(27 downto 0); 
            SV41_dim5 : in std_logic_vector(27 downto 0); 
            SV41_dim6 : in std_logic_vector(27 downto 0); 
            SV41_dim7 : in std_logic_vector(27 downto 0); 
            SV42_dim0 : in std_logic_vector(27 downto 0); 
            SV42_dim1 : in std_logic_vector(27 downto 0); 
            SV42_dim2 : in std_logic_vector(27 downto 0); 
            SV42_dim3 : in std_logic_vector(27 downto 0); 
            SV42_dim4 : in std_logic_vector(27 downto 0); 
            SV42_dim5 : in std_logic_vector(27 downto 0); 
            SV42_dim6 : in std_logic_vector(27 downto 0); 
            SV42_dim7 : in std_logic_vector(27 downto 0); 
            SV43_dim0 : in std_logic_vector(27 downto 0); 
            SV43_dim1 : in std_logic_vector(27 downto 0); 
            SV43_dim2 : in std_logic_vector(27 downto 0); 
            SV43_dim3 : in std_logic_vector(27 downto 0); 
            SV43_dim4 : in std_logic_vector(27 downto 0); 
            SV43_dim5 : in std_logic_vector(27 downto 0); 
            SV43_dim6 : in std_logic_vector(27 downto 0); 
            SV43_dim7 : in std_logic_vector(27 downto 0); 
            SV44_dim0 : in std_logic_vector(27 downto 0); 
            SV44_dim1 : in std_logic_vector(27 downto 0); 
            SV44_dim2 : in std_logic_vector(27 downto 0); 
            SV44_dim3 : in std_logic_vector(27 downto 0); 
            SV44_dim4 : in std_logic_vector(27 downto 0); 
            SV44_dim5 : in std_logic_vector(27 downto 0); 
            SV44_dim6 : in std_logic_vector(27 downto 0); 
            SV44_dim7 : in std_logic_vector(27 downto 0); 
            SV45_dim0 : in std_logic_vector(27 downto 0); 
            SV45_dim1 : in std_logic_vector(27 downto 0); 
            SV45_dim2 : in std_logic_vector(27 downto 0); 
            SV45_dim3 : in std_logic_vector(27 downto 0); 
            SV45_dim4 : in std_logic_vector(27 downto 0); 
            SV45_dim5 : in std_logic_vector(27 downto 0); 
            SV45_dim6 : in std_logic_vector(27 downto 0); 
            SV45_dim7 : in std_logic_vector(27 downto 0); 
            SV46_dim0 : in std_logic_vector(27 downto 0); 
            SV46_dim1 : in std_logic_vector(27 downto 0); 
            SV46_dim2 : in std_logic_vector(27 downto 0); 
            SV46_dim3 : in std_logic_vector(27 downto 0); 
            SV46_dim4 : in std_logic_vector(27 downto 0); 
            SV46_dim5 : in std_logic_vector(27 downto 0); 
            SV46_dim6 : in std_logic_vector(27 downto 0); 
            SV46_dim7 : in std_logic_vector(27 downto 0); 
            SV47_dim0 : in std_logic_vector(27 downto 0); 
            SV47_dim1 : in std_logic_vector(27 downto 0); 
            SV47_dim2 : in std_logic_vector(27 downto 0); 
            SV47_dim3 : in std_logic_vector(27 downto 0); 
            SV47_dim4 : in std_logic_vector(27 downto 0); 
            SV47_dim5 : in std_logic_vector(27 downto 0); 
            SV47_dim6 : in std_logic_vector(27 downto 0); 
            SV47_dim7 : in std_logic_vector(27 downto 0); 
            SV48_dim0 : in std_logic_vector(27 downto 0); 
            SV48_dim1 : in std_logic_vector(27 downto 0); 
            SV48_dim2 : in std_logic_vector(27 downto 0); 
            SV48_dim3 : in std_logic_vector(27 downto 0); 
            SV48_dim4 : in std_logic_vector(27 downto 0); 
            SV48_dim5 : in std_logic_vector(27 downto 0); 
            SV48_dim6 : in std_logic_vector(27 downto 0); 
            SV48_dim7 : in std_logic_vector(27 downto 0); 
            SV49_dim0 : in std_logic_vector(27 downto 0); 
            SV49_dim1 : in std_logic_vector(27 downto 0); 
            SV49_dim2 : in std_logic_vector(27 downto 0); 
            SV49_dim3 : in std_logic_vector(27 downto 0); 
            SV49_dim4 : in std_logic_vector(27 downto 0); 
            SV49_dim5 : in std_logic_vector(27 downto 0); 
            SV49_dim6 : in std_logic_vector(27 downto 0); 
            SV49_dim7 : in std_logic_vector(27 downto 0); 
            SV50_dim0 : in std_logic_vector(27 downto 0); 
            SV50_dim1 : in std_logic_vector(27 downto 0); 
            SV50_dim2 : in std_logic_vector(27 downto 0); 
            SV50_dim3 : in std_logic_vector(27 downto 0); 
            SV50_dim4 : in std_logic_vector(27 downto 0); 
            SV50_dim5 : in std_logic_vector(27 downto 0); 
            SV50_dim6 : in std_logic_vector(27 downto 0); 
            SV50_dim7 : in std_logic_vector(27 downto 0); 
            SV51_dim0 : in std_logic_vector(27 downto 0); 
            SV51_dim1 : in std_logic_vector(27 downto 0); 
            SV51_dim2 : in std_logic_vector(27 downto 0); 
            SV51_dim3 : in std_logic_vector(27 downto 0); 
            SV51_dim4 : in std_logic_vector(27 downto 0); 
            SV51_dim5 : in std_logic_vector(27 downto 0); 
            SV51_dim6 : in std_logic_vector(27 downto 0); 
            SV51_dim7 : in std_logic_vector(27 downto 0); 
            SV52_dim0 : in std_logic_vector(27 downto 0); 
            SV52_dim1 : in std_logic_vector(27 downto 0); 
            SV52_dim2 : in std_logic_vector(27 downto 0); 
            SV52_dim3 : in std_logic_vector(27 downto 0); 
            SV52_dim4 : in std_logic_vector(27 downto 0); 
            SV52_dim5 : in std_logic_vector(27 downto 0); 
            SV52_dim6 : in std_logic_vector(27 downto 0); 
            SV52_dim7 : in std_logic_vector(27 downto 0); 
            SV53_dim0 : in std_logic_vector(27 downto 0); 
            SV53_dim1 : in std_logic_vector(27 downto 0); 
            SV53_dim2 : in std_logic_vector(27 downto 0); 
            SV53_dim3 : in std_logic_vector(27 downto 0); 
            SV53_dim4 : in std_logic_vector(27 downto 0); 
            SV53_dim5 : in std_logic_vector(27 downto 0); 
            SV53_dim6 : in std_logic_vector(27 downto 0); 
            SV53_dim7 : in std_logic_vector(27 downto 0); 
            SV54_dim0 : in std_logic_vector(27 downto 0); 
            SV54_dim1 : in std_logic_vector(27 downto 0); 
            SV54_dim2 : in std_logic_vector(27 downto 0); 
            SV54_dim3 : in std_logic_vector(27 downto 0); 
            SV54_dim4 : in std_logic_vector(27 downto 0); 
            SV54_dim5 : in std_logic_vector(27 downto 0); 
            SV54_dim6 : in std_logic_vector(27 downto 0); 
            SV54_dim7 : in std_logic_vector(27 downto 0); 
            SV55_dim0 : in std_logic_vector(27 downto 0); 
            SV55_dim1 : in std_logic_vector(27 downto 0); 
            SV55_dim2 : in std_logic_vector(27 downto 0); 
            SV55_dim3 : in std_logic_vector(27 downto 0); 
            SV55_dim4 : in std_logic_vector(27 downto 0); 
            SV55_dim5 : in std_logic_vector(27 downto 0); 
            SV55_dim6 : in std_logic_vector(27 downto 0); 
            SV55_dim7 : in std_logic_vector(27 downto 0); 
            SV56_dim0 : in std_logic_vector(27 downto 0); 
            SV56_dim1 : in std_logic_vector(27 downto 0); 
            SV56_dim2 : in std_logic_vector(27 downto 0); 
            SV56_dim3 : in std_logic_vector(27 downto 0); 
            SV56_dim4 : in std_logic_vector(27 downto 0); 
            SV56_dim5 : in std_logic_vector(27 downto 0); 
            SV56_dim6 : in std_logic_vector(27 downto 0); 
            SV56_dim7 : in std_logic_vector(27 downto 0); 
            SV57_dim0 : in std_logic_vector(27 downto 0); 
            SV57_dim1 : in std_logic_vector(27 downto 0); 
            SV57_dim2 : in std_logic_vector(27 downto 0); 
            SV57_dim3 : in std_logic_vector(27 downto 0); 
            SV57_dim4 : in std_logic_vector(27 downto 0); 
            SV57_dim5 : in std_logic_vector(27 downto 0); 
            SV57_dim6 : in std_logic_vector(27 downto 0); 
            SV57_dim7 : in std_logic_vector(27 downto 0); 
            SV58_dim0 : in std_logic_vector(27 downto 0); 
            SV58_dim1 : in std_logic_vector(27 downto 0); 
            SV58_dim2 : in std_logic_vector(27 downto 0); 
            SV58_dim3 : in std_logic_vector(27 downto 0); 
            SV58_dim4 : in std_logic_vector(27 downto 0); 
            SV58_dim5 : in std_logic_vector(27 downto 0); 
            SV58_dim6 : in std_logic_vector(27 downto 0); 
            SV58_dim7 : in std_logic_vector(27 downto 0); 
            SV59_dim0 : in std_logic_vector(27 downto 0); 
            SV59_dim1 : in std_logic_vector(27 downto 0); 
            SV59_dim2 : in std_logic_vector(27 downto 0); 
            SV59_dim3 : in std_logic_vector(27 downto 0); 
            SV59_dim4 : in std_logic_vector(27 downto 0); 
            SV59_dim5 : in std_logic_vector(27 downto 0); 
            SV59_dim6 : in std_logic_vector(27 downto 0); 
            SV59_dim7 : in std_logic_vector(27 downto 0); 
            SV60_dim0 : in std_logic_vector(27 downto 0); 
            SV60_dim1 : in std_logic_vector(27 downto 0); 
            SV60_dim2 : in std_logic_vector(27 downto 0); 
            SV60_dim3 : in std_logic_vector(27 downto 0); 
            SV60_dim4 : in std_logic_vector(27 downto 0); 
            SV60_dim5 : in std_logic_vector(27 downto 0); 
            SV60_dim6 : in std_logic_vector(27 downto 0); 
            SV60_dim7 : in std_logic_vector(27 downto 0); 
            SV61_dim0 : in std_logic_vector(27 downto 0); 
            SV61_dim1 : in std_logic_vector(27 downto 0); 
            SV61_dim2 : in std_logic_vector(27 downto 0); 
            SV61_dim3 : in std_logic_vector(27 downto 0); 
            SV61_dim4 : in std_logic_vector(27 downto 0); 
            SV61_dim5 : in std_logic_vector(27 downto 0); 
            SV61_dim6 : in std_logic_vector(27 downto 0); 
            SV61_dim7 : in std_logic_vector(27 downto 0); 
            SV62_dim0 : in std_logic_vector(27 downto 0); 
            SV62_dim1 : in std_logic_vector(27 downto 0); 
            SV62_dim2 : in std_logic_vector(27 downto 0); 
            SV62_dim3 : in std_logic_vector(27 downto 0); 
            SV62_dim4 : in std_logic_vector(27 downto 0); 
            SV62_dim5 : in std_logic_vector(27 downto 0); 
            SV62_dim6 : in std_logic_vector(27 downto 0); 
            SV62_dim7 : in std_logic_vector(27 downto 0); 
            SV63_dim0 : in std_logic_vector(27 downto 0); 
            SV63_dim1 : in std_logic_vector(27 downto 0); 
            SV63_dim2 : in std_logic_vector(27 downto 0); 
            SV63_dim3 : in std_logic_vector(27 downto 0); 
            SV63_dim4 : in std_logic_vector(27 downto 0); 
            SV63_dim5 : in std_logic_vector(27 downto 0); 
            SV63_dim6 : in std_logic_vector(27 downto 0); 
            SV63_dim7 : in std_logic_vector(27 downto 0); 
            SV64_dim0 : in std_logic_vector(27 downto 0); 
            SV64_dim1 : in std_logic_vector(27 downto 0); 
            SV64_dim2 : in std_logic_vector(27 downto 0); 
            SV64_dim3 : in std_logic_vector(27 downto 0); 
            SV64_dim4 : in std_logic_vector(27 downto 0); 
            SV64_dim5 : in std_logic_vector(27 downto 0); 
            SV64_dim6 : in std_logic_vector(27 downto 0); 
            SV64_dim7 : in std_logic_vector(27 downto 0); 
            SV65_dim0 : in std_logic_vector(27 downto 0); 
            SV65_dim1 : in std_logic_vector(27 downto 0); 
            SV65_dim2 : in std_logic_vector(27 downto 0); 
            SV65_dim3 : in std_logic_vector(27 downto 0); 
            SV65_dim4 : in std_logic_vector(27 downto 0); 
            SV65_dim5 : in std_logic_vector(27 downto 0); 
            SV65_dim6 : in std_logic_vector(27 downto 0); 
            SV65_dim7 : in std_logic_vector(27 downto 0); 
            SV66_dim0 : in std_logic_vector(27 downto 0); 
            SV66_dim1 : in std_logic_vector(27 downto 0); 
            SV66_dim2 : in std_logic_vector(27 downto 0); 
            SV66_dim3 : in std_logic_vector(27 downto 0); 
            SV66_dim4 : in std_logic_vector(27 downto 0); 
            SV66_dim5 : in std_logic_vector(27 downto 0); 
            SV66_dim6 : in std_logic_vector(27 downto 0); 
            SV66_dim7 : in std_logic_vector(27 downto 0); 
            SV67_dim0 : in std_logic_vector(27 downto 0); 
            SV67_dim1 : in std_logic_vector(27 downto 0); 
            SV67_dim2 : in std_logic_vector(27 downto 0); 
            SV67_dim3 : in std_logic_vector(27 downto 0); 
            SV67_dim4 : in std_logic_vector(27 downto 0); 
            SV67_dim5 : in std_logic_vector(27 downto 0); 
            SV67_dim6 : in std_logic_vector(27 downto 0); 
            SV67_dim7 : in std_logic_vector(27 downto 0); 
            SV68_dim0 : in std_logic_vector(27 downto 0); 
            SV68_dim1 : in std_logic_vector(27 downto 0); 
            SV68_dim2 : in std_logic_vector(27 downto 0); 
            SV68_dim3 : in std_logic_vector(27 downto 0); 
            SV68_dim4 : in std_logic_vector(27 downto 0); 
            SV68_dim5 : in std_logic_vector(27 downto 0); 
            SV68_dim6 : in std_logic_vector(27 downto 0); 
            SV68_dim7 : in std_logic_vector(27 downto 0); 
            SV69_dim0 : in std_logic_vector(27 downto 0); 
            SV69_dim1 : in std_logic_vector(27 downto 0); 
            SV69_dim2 : in std_logic_vector(27 downto 0); 
            SV69_dim3 : in std_logic_vector(27 downto 0); 
            SV69_dim4 : in std_logic_vector(27 downto 0); 
            SV69_dim5 : in std_logic_vector(27 downto 0); 
            SV69_dim6 : in std_logic_vector(27 downto 0); 
            SV69_dim7 : in std_logic_vector(27 downto 0); 
            SV70_dim0 : in std_logic_vector(27 downto 0); 
            SV70_dim1 : in std_logic_vector(27 downto 0); 
            SV70_dim2 : in std_logic_vector(27 downto 0); 
            SV70_dim3 : in std_logic_vector(27 downto 0); 
            SV70_dim4 : in std_logic_vector(27 downto 0); 
            SV70_dim5 : in std_logic_vector(27 downto 0); 
            SV70_dim6 : in std_logic_vector(27 downto 0); 
            SV70_dim7 : in std_logic_vector(27 downto 0); 
            
            -- Test Data
            test_data_dim0 : in std_logic_vector(27 downto 0); 
            test_data_dim1 : in std_logic_vector(27 downto 0); 
            test_data_dim2 : in std_logic_vector(27 downto 0); 
            test_data_dim3 : in std_logic_vector(27 downto 0); 
            test_data_dim4 : in std_logic_vector(27 downto 0); 
            test_data_dim5 : in std_logic_vector(27 downto 0); 
            test_data_dim6 : in std_logic_vector(27 downto 0); 
            test_data_dim7 : in std_logic_vector(27 downto 0); 
            
            -- alpha * Y
			SV0_alphaY : in std_logic_vector(11 downto 0); 
			SV1_alphaY : in std_logic_vector(11 downto 0); 
			SV2_alphaY : in std_logic_vector(11 downto 0); 
			SV3_alphaY : in std_logic_vector(11 downto 0); 
			SV4_alphaY : in std_logic_vector(11 downto 0); 
			SV5_alphaY : in std_logic_vector(11 downto 0); 
			SV6_alphaY : in std_logic_vector(11 downto 0); 
			SV7_alphaY : in std_logic_vector(11 downto 0); 
			SV8_alphaY : in std_logic_vector(11 downto 0); 
			SV9_alphaY : in std_logic_vector(11 downto 0); 
			SV10_alphaY : in std_logic_vector(11 downto 0); 
			SV11_alphaY : in std_logic_vector(11 downto 0); 
			SV12_alphaY : in std_logic_vector(11 downto 0); 
			SV13_alphaY : in std_logic_vector(11 downto 0); 
			SV14_alphaY : in std_logic_vector(11 downto 0); 
			SV15_alphaY : in std_logic_vector(11 downto 0); 
			SV16_alphaY : in std_logic_vector(11 downto 0); 
			SV17_alphaY : in std_logic_vector(11 downto 0); 
			SV18_alphaY : in std_logic_vector(11 downto 0); 
			SV19_alphaY : in std_logic_vector(11 downto 0); 
			SV20_alphaY : in std_logic_vector(11 downto 0); 
			SV21_alphaY : in std_logic_vector(11 downto 0); 
			SV22_alphaY : in std_logic_vector(11 downto 0); 
			SV23_alphaY : in std_logic_vector(11 downto 0); 
			SV24_alphaY : in std_logic_vector(11 downto 0); 
			SV25_alphaY : in std_logic_vector(11 downto 0); 
			SV26_alphaY : in std_logic_vector(11 downto 0); 
			SV27_alphaY : in std_logic_vector(11 downto 0); 
			SV28_alphaY : in std_logic_vector(11 downto 0); 
			SV29_alphaY : in std_logic_vector(11 downto 0); 
			SV30_alphaY : in std_logic_vector(11 downto 0); 
			SV31_alphaY : in std_logic_vector(11 downto 0); 
			SV32_alphaY : in std_logic_vector(11 downto 0); 
			SV33_alphaY : in std_logic_vector(11 downto 0); 
			SV34_alphaY : in std_logic_vector(11 downto 0); 
			SV35_alphaY : in std_logic_vector(11 downto 0); 
			SV36_alphaY : in std_logic_vector(11 downto 0); 
			SV37_alphaY : in std_logic_vector(11 downto 0); 
			SV38_alphaY : in std_logic_vector(11 downto 0); 
			SV39_alphaY : in std_logic_vector(11 downto 0); 
			SV40_alphaY : in std_logic_vector(11 downto 0); 
			SV41_alphaY : in std_logic_vector(11 downto 0); 
			SV42_alphaY : in std_logic_vector(11 downto 0); 
			SV43_alphaY : in std_logic_vector(11 downto 0); 
			SV44_alphaY : in std_logic_vector(11 downto 0); 
			SV45_alphaY : in std_logic_vector(11 downto 0); 
			SV46_alphaY : in std_logic_vector(11 downto 0); 
			SV47_alphaY : in std_logic_vector(11 downto 0); 
			SV48_alphaY : in std_logic_vector(11 downto 0); 
			SV49_alphaY : in std_logic_vector(11 downto 0); 
			SV50_alphaY : in std_logic_vector(11 downto 0); 
			SV51_alphaY : in std_logic_vector(11 downto 0); 
			SV52_alphaY : in std_logic_vector(11 downto 0); 
			SV53_alphaY : in std_logic_vector(11 downto 0); 
			SV54_alphaY : in std_logic_vector(11 downto 0); 
			SV55_alphaY : in std_logic_vector(11 downto 0); 
			SV56_alphaY : in std_logic_vector(11 downto 0); 
			SV57_alphaY : in std_logic_vector(11 downto 0); 
			SV58_alphaY : in std_logic_vector(11 downto 0); 
			SV59_alphaY : in std_logic_vector(11 downto 0); 
			SV60_alphaY : in std_logic_vector(11 downto 0); 
			SV61_alphaY : in std_logic_vector(11 downto 0); 
			SV62_alphaY : in std_logic_vector(11 downto 0); 
			SV63_alphaY : in std_logic_vector(11 downto 0); 
			SV64_alphaY : in std_logic_vector(11 downto 0); 
			SV65_alphaY : in std_logic_vector(11 downto 0); 
			SV66_alphaY : in std_logic_vector(11 downto 0); 
			SV67_alphaY : in std_logic_vector(11 downto 0); 
			SV68_alphaY : in std_logic_vector(11 downto 0); 
			SV69_alphaY : in std_logic_vector(11 downto 0); 
			SV70_alphaY : in std_logic_vector(11 downto 0); 
            
            -- gamma
            gamma : in std_logic_vector(11 downto 0); 
            
            -- b
            b : in std_logic_vector(19 downto 0); 
            
            -- output
            output : out std_logic
            );
end TOP;

architecture Behavioral of TOP is

component Kernel_rbf is
    Port (  SV_dim0 : in std_logic_vector(27 downto 0);
            SV_dim1 : in std_logic_vector(27 downto 0);
            SV_dim2 : in std_logic_vector(27 downto 0);
            SV_dim3 : in std_logic_vector(27 downto 0);
            SV_dim4 : in std_logic_vector(27 downto 0);
            SV_dim5 : in std_logic_vector(27 downto 0);
            SV_dim6 : in std_logic_vector(27 downto 0);
            SV_dim7 : in std_logic_vector(27 downto 0);
            test_data_dim0 : in std_logic_vector(27 downto 0);
            test_data_dim1 : in std_logic_vector(27 downto 0);
            test_data_dim2 : in std_logic_vector(27 downto 0);
            test_data_dim3 : in std_logic_vector(27 downto 0);
            test_data_dim4 : in std_logic_vector(27 downto 0);
            test_data_dim5 : in std_logic_vector(27 downto 0);
            test_data_dim6 : in std_logic_vector(27 downto 0);
            test_data_dim7 : in std_logic_vector(27 downto 0);
            gamma : in std_logic_vector(11 downto 0);
            output : out std_logic_vector(10 downto 0)
            );
end component;

component Multiplier_Signed_12bits is
    Port (  input_a : in std_logic_vector(11 downto 0);     
            input_b : in std_logic_vector(11 downto 0);
            output : out std_logic_vector(12 downto 0)  -- (SIGNED)2bit.10bits * (SIGNED)2bit.10bits = (SIGNED)3bits.10bits
            );
end component;

component Adder_Signed_20bits is
    Port (  input_a : in std_logic_vector(19 downto 0);
            input_b : in std_logic_vector(19 downto 0);
            output : out std_logic_vector(19 downto 0);
            overflow : out std_logic
            );
end component;

-- Kernel_rbf Signal
signal Kernel_rbf_output_s0 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s1 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s2 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s3 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s4 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s5 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s6 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s7 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s8 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s9 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s10 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s11 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s12 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s13 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s14 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s15 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s16 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s17 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s18 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s19 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s20 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s21 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s22 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s23 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s24 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s25 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s26 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s27 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s28 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s29 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s30 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s31 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s32 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s33 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s34 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s35 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s36 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s37 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s38 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s39 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s40 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s41 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s42 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s43 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s44 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s45 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s46 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s47 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s48 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s49 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s50 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s51 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s52 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s53 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s54 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s55 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s56 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s57 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s58 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s59 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s60 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s61 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s62 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s63 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s64 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s65 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s66 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s67 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s68 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s69 : std_logic_vector(10 downto 0); 
signal Kernel_rbf_output_s70 : std_logic_vector(10 downto 0); 

-- Multiplier Signal
signal multi_s0 : std_logic_vector(12 downto 0);
signal multi_s1 : std_logic_vector(12 downto 0);
signal multi_s2 : std_logic_vector(12 downto 0);
signal multi_s3 : std_logic_vector(12 downto 0);
signal multi_s4 : std_logic_vector(12 downto 0);
signal multi_s5 : std_logic_vector(12 downto 0);
signal multi_s6 : std_logic_vector(12 downto 0);
signal multi_s7 : std_logic_vector(12 downto 0);
signal multi_s8 : std_logic_vector(12 downto 0);
signal multi_s9 : std_logic_vector(12 downto 0);
signal multi_s10 : std_logic_vector(12 downto 0);
signal multi_s11 : std_logic_vector(12 downto 0);
signal multi_s12 : std_logic_vector(12 downto 0);
signal multi_s13 : std_logic_vector(12 downto 0);
signal multi_s14 : std_logic_vector(12 downto 0);
signal multi_s15 : std_logic_vector(12 downto 0);
signal multi_s16 : std_logic_vector(12 downto 0);
signal multi_s17 : std_logic_vector(12 downto 0);
signal multi_s18 : std_logic_vector(12 downto 0);
signal multi_s19 : std_logic_vector(12 downto 0);
signal multi_s20 : std_logic_vector(12 downto 0);
signal multi_s21 : std_logic_vector(12 downto 0);
signal multi_s22 : std_logic_vector(12 downto 0);
signal multi_s23 : std_logic_vector(12 downto 0);
signal multi_s24 : std_logic_vector(12 downto 0);
signal multi_s25 : std_logic_vector(12 downto 0);
signal multi_s26 : std_logic_vector(12 downto 0);
signal multi_s27 : std_logic_vector(12 downto 0);
signal multi_s28 : std_logic_vector(12 downto 0);
signal multi_s29 : std_logic_vector(12 downto 0);
signal multi_s30 : std_logic_vector(12 downto 0);
signal multi_s31 : std_logic_vector(12 downto 0);
signal multi_s32 : std_logic_vector(12 downto 0);
signal multi_s33 : std_logic_vector(12 downto 0);
signal multi_s34 : std_logic_vector(12 downto 0);
signal multi_s35 : std_logic_vector(12 downto 0);
signal multi_s36 : std_logic_vector(12 downto 0);
signal multi_s37 : std_logic_vector(12 downto 0);
signal multi_s38 : std_logic_vector(12 downto 0);
signal multi_s39 : std_logic_vector(12 downto 0);
signal multi_s40 : std_logic_vector(12 downto 0);
signal multi_s41 : std_logic_vector(12 downto 0);
signal multi_s42 : std_logic_vector(12 downto 0);
signal multi_s43 : std_logic_vector(12 downto 0);
signal multi_s44 : std_logic_vector(12 downto 0);
signal multi_s45 : std_logic_vector(12 downto 0);
signal multi_s46 : std_logic_vector(12 downto 0);
signal multi_s47 : std_logic_vector(12 downto 0);
signal multi_s48 : std_logic_vector(12 downto 0);
signal multi_s49 : std_logic_vector(12 downto 0);
signal multi_s50 : std_logic_vector(12 downto 0);
signal multi_s51 : std_logic_vector(12 downto 0);
signal multi_s52 : std_logic_vector(12 downto 0);
signal multi_s53 : std_logic_vector(12 downto 0);
signal multi_s54 : std_logic_vector(12 downto 0);
signal multi_s55 : std_logic_vector(12 downto 0);
signal multi_s56 : std_logic_vector(12 downto 0);
signal multi_s57 : std_logic_vector(12 downto 0);
signal multi_s58 : std_logic_vector(12 downto 0);
signal multi_s59 : std_logic_vector(12 downto 0);
signal multi_s60 : std_logic_vector(12 downto 0);
signal multi_s61 : std_logic_vector(12 downto 0);
signal multi_s62 : std_logic_vector(12 downto 0);
signal multi_s63 : std_logic_vector(12 downto 0);
signal multi_s64 : std_logic_vector(12 downto 0);
signal multi_s65 : std_logic_vector(12 downto 0);
signal multi_s66 : std_logic_vector(12 downto 0);
signal multi_s67 : std_logic_vector(12 downto 0);
signal multi_s68 : std_logic_vector(12 downto 0);
signal multi_s69 : std_logic_vector(12 downto 0);
signal multi_s70 : std_logic_vector(12 downto 0);

-- Adder Signal
signal add_output_s00 : std_logic_vector(19 downto 0); 
signal add_output_s01 : std_logic_vector(19 downto 0); 
signal add_output_s02 : std_logic_vector(19 downto 0); 
signal add_output_s03 : std_logic_vector(19 downto 0); 
signal add_output_s04 : std_logic_vector(19 downto 0); 
signal add_output_s05 : std_logic_vector(19 downto 0); 
signal add_output_s06 : std_logic_vector(19 downto 0); 
signal add_output_s07 : std_logic_vector(19 downto 0); 
signal add_output_s08 : std_logic_vector(19 downto 0); 
signal add_output_s09 : std_logic_vector(19 downto 0); 
signal add_output_s010 : std_logic_vector(19 downto 0); 
signal add_output_s011 : std_logic_vector(19 downto 0); 
signal add_output_s012 : std_logic_vector(19 downto 0); 
signal add_output_s013 : std_logic_vector(19 downto 0); 
signal add_output_s014 : std_logic_vector(19 downto 0); 
signal add_output_s015 : std_logic_vector(19 downto 0); 
signal add_output_s016 : std_logic_vector(19 downto 0); 
signal add_output_s017 : std_logic_vector(19 downto 0); 
signal add_output_s018 : std_logic_vector(19 downto 0); 
signal add_output_s019 : std_logic_vector(19 downto 0); 
signal add_output_s020 : std_logic_vector(19 downto 0); 
signal add_output_s021 : std_logic_vector(19 downto 0); 
signal add_output_s022 : std_logic_vector(19 downto 0); 
signal add_output_s023 : std_logic_vector(19 downto 0); 
signal add_output_s024 : std_logic_vector(19 downto 0); 
signal add_output_s025 : std_logic_vector(19 downto 0); 
signal add_output_s026 : std_logic_vector(19 downto 0); 
signal add_output_s027 : std_logic_vector(19 downto 0); 
signal add_output_s028 : std_logic_vector(19 downto 0); 
signal add_output_s029 : std_logic_vector(19 downto 0); 
signal add_output_s030 : std_logic_vector(19 downto 0); 
signal add_output_s031 : std_logic_vector(19 downto 0); 
signal add_output_s032 : std_logic_vector(19 downto 0); 
signal add_output_s033 : std_logic_vector(19 downto 0); 
signal add_output_s034 : std_logic_vector(19 downto 0); 
signal add_output_s035 : std_logic_vector(19 downto 0); 
signal add_output_s10 : std_logic_vector(19 downto 0); 
signal add_output_s11 : std_logic_vector(19 downto 0); 
signal add_output_s12 : std_logic_vector(19 downto 0); 
signal add_output_s13 : std_logic_vector(19 downto 0); 
signal add_output_s14 : std_logic_vector(19 downto 0); 
signal add_output_s15 : std_logic_vector(19 downto 0); 
signal add_output_s16 : std_logic_vector(19 downto 0); 
signal add_output_s17 : std_logic_vector(19 downto 0); 
signal add_output_s18 : std_logic_vector(19 downto 0); 
signal add_output_s19 : std_logic_vector(19 downto 0); 
signal add_output_s110 : std_logic_vector(19 downto 0); 
signal add_output_s111 : std_logic_vector(19 downto 0); 
signal add_output_s112 : std_logic_vector(19 downto 0); 
signal add_output_s113 : std_logic_vector(19 downto 0); 
signal add_output_s114 : std_logic_vector(19 downto 0); 
signal add_output_s115 : std_logic_vector(19 downto 0); 
signal add_output_s116 : std_logic_vector(19 downto 0); 
signal add_output_s117 : std_logic_vector(19 downto 0); 
signal add_output_s20 : std_logic_vector(19 downto 0); 
signal add_output_s21 : std_logic_vector(19 downto 0); 
signal add_output_s22 : std_logic_vector(19 downto 0); 
signal add_output_s23 : std_logic_vector(19 downto 0); 
signal add_output_s24 : std_logic_vector(19 downto 0); 
signal add_output_s25 : std_logic_vector(19 downto 0); 
signal add_output_s26 : std_logic_vector(19 downto 0); 
signal add_output_s27 : std_logic_vector(19 downto 0); 
signal add_output_s28 : std_logic_vector(19 downto 0); 
signal add_output_s30 : std_logic_vector(19 downto 0); 
signal add_output_s31 : std_logic_vector(19 downto 0); 
signal add_output_s32 : std_logic_vector(19 downto 0); 
signal add_output_s33 : std_logic_vector(19 downto 0); 
signal add_output_s40 : std_logic_vector(19 downto 0); 
signal add_output_s41 : std_logic_vector(19 downto 0); 
signal add_output_s50 : std_logic_vector(19 downto 0); 
signal add_output_s60 : std_logic_vector(19 downto 0); 
signal add_overflow_s00 : std_logic; 
signal add_overflow_s01 : std_logic; 
signal add_overflow_s02 : std_logic; 
signal add_overflow_s03 : std_logic; 
signal add_overflow_s04 : std_logic; 
signal add_overflow_s05 : std_logic; 
signal add_overflow_s06 : std_logic; 
signal add_overflow_s07 : std_logic; 
signal add_overflow_s08 : std_logic; 
signal add_overflow_s09 : std_logic; 
signal add_overflow_s010 : std_logic; 
signal add_overflow_s011 : std_logic; 
signal add_overflow_s012 : std_logic; 
signal add_overflow_s013 : std_logic; 
signal add_overflow_s014 : std_logic; 
signal add_overflow_s015 : std_logic; 
signal add_overflow_s016 : std_logic; 
signal add_overflow_s017 : std_logic; 
signal add_overflow_s018 : std_logic; 
signal add_overflow_s019 : std_logic; 
signal add_overflow_s020 : std_logic; 
signal add_overflow_s021 : std_logic; 
signal add_overflow_s022 : std_logic; 
signal add_overflow_s023 : std_logic; 
signal add_overflow_s024 : std_logic; 
signal add_overflow_s025 : std_logic; 
signal add_overflow_s026 : std_logic; 
signal add_overflow_s027 : std_logic; 
signal add_overflow_s028 : std_logic; 
signal add_overflow_s029 : std_logic; 
signal add_overflow_s030 : std_logic; 
signal add_overflow_s031 : std_logic; 
signal add_overflow_s032 : std_logic; 
signal add_overflow_s033 : std_logic; 
signal add_overflow_s034 : std_logic; 
signal add_overflow_s035 : std_logic; 
signal add_overflow_s10 : std_logic; 
signal add_overflow_s11 : std_logic; 
signal add_overflow_s12 : std_logic; 
signal add_overflow_s13 : std_logic; 
signal add_overflow_s14 : std_logic; 
signal add_overflow_s15 : std_logic; 
signal add_overflow_s16 : std_logic; 
signal add_overflow_s17 : std_logic; 
signal add_overflow_s18 : std_logic; 
signal add_overflow_s19 : std_logic; 
signal add_overflow_s110 : std_logic; 
signal add_overflow_s111 : std_logic; 
signal add_overflow_s112 : std_logic; 
signal add_overflow_s113 : std_logic; 
signal add_overflow_s114 : std_logic; 
signal add_overflow_s115 : std_logic; 
signal add_overflow_s116 : std_logic; 
signal add_overflow_s117 : std_logic; 
signal add_overflow_s20 : std_logic; 
signal add_overflow_s21 : std_logic; 
signal add_overflow_s22 : std_logic; 
signal add_overflow_s23 : std_logic; 
signal add_overflow_s24 : std_logic; 
signal add_overflow_s25 : std_logic; 
signal add_overflow_s26 : std_logic; 
signal add_overflow_s27 : std_logic; 
signal add_overflow_s28 : std_logic; 
signal add_overflow_s30 : std_logic; 
signal add_overflow_s31 : std_logic; 
signal add_overflow_s32 : std_logic; 
signal add_overflow_s33 : std_logic; 
signal add_overflow_s40 : std_logic; 
signal add_overflow_s41 : std_logic; 
signal add_overflow_s50 : std_logic; 
signal add_overflow_s60 : std_logic;     

begin

	Kernel_rbf_0 : Kernel_rbf
	port map(	SV_dim0 => SV0_dim0,
				SV_dim1 => SV0_dim1,
				SV_dim2 => SV0_dim2,
				SV_dim3 => SV0_dim3,
				SV_dim4 => SV0_dim4,
				SV_dim5 => SV0_dim5,
				SV_dim6 => SV0_dim6,
				SV_dim7 => SV0_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s0
				);

	Kernel_rbf_1 : Kernel_rbf
	port map(	SV_dim0 => SV1_dim0,
				SV_dim1 => SV1_dim1,
				SV_dim2 => SV1_dim2,
				SV_dim3 => SV1_dim3,
				SV_dim4 => SV1_dim4,
				SV_dim5 => SV1_dim5,
				SV_dim6 => SV1_dim6,
				SV_dim7 => SV1_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s1
				);

	Kernel_rbf_2 : Kernel_rbf
	port map(	SV_dim0 => SV2_dim0,
				SV_dim1 => SV2_dim1,
				SV_dim2 => SV2_dim2,
				SV_dim3 => SV2_dim3,
				SV_dim4 => SV2_dim4,
				SV_dim5 => SV2_dim5,
				SV_dim6 => SV2_dim6,
				SV_dim7 => SV2_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s2
				);

	Kernel_rbf_3 : Kernel_rbf
	port map(	SV_dim0 => SV3_dim0,
				SV_dim1 => SV3_dim1,
				SV_dim2 => SV3_dim2,
				SV_dim3 => SV3_dim3,
				SV_dim4 => SV3_dim4,
				SV_dim5 => SV3_dim5,
				SV_dim6 => SV3_dim6,
				SV_dim7 => SV3_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s3
				);

	Kernel_rbf_4 : Kernel_rbf
	port map(	SV_dim0 => SV4_dim0,
				SV_dim1 => SV4_dim1,
				SV_dim2 => SV4_dim2,
				SV_dim3 => SV4_dim3,
				SV_dim4 => SV4_dim4,
				SV_dim5 => SV4_dim5,
				SV_dim6 => SV4_dim6,
				SV_dim7 => SV4_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s4
				);

	Kernel_rbf_5 : Kernel_rbf
	port map(	SV_dim0 => SV5_dim0,
				SV_dim1 => SV5_dim1,
				SV_dim2 => SV5_dim2,
				SV_dim3 => SV5_dim3,
				SV_dim4 => SV5_dim4,
				SV_dim5 => SV5_dim5,
				SV_dim6 => SV5_dim6,
				SV_dim7 => SV5_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s5
				);

	Kernel_rbf_6 : Kernel_rbf
	port map(	SV_dim0 => SV6_dim0,
				SV_dim1 => SV6_dim1,
				SV_dim2 => SV6_dim2,
				SV_dim3 => SV6_dim3,
				SV_dim4 => SV6_dim4,
				SV_dim5 => SV6_dim5,
				SV_dim6 => SV6_dim6,
				SV_dim7 => SV6_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s6
				);

	Kernel_rbf_7 : Kernel_rbf
	port map(	SV_dim0 => SV7_dim0,
				SV_dim1 => SV7_dim1,
				SV_dim2 => SV7_dim2,
				SV_dim3 => SV7_dim3,
				SV_dim4 => SV7_dim4,
				SV_dim5 => SV7_dim5,
				SV_dim6 => SV7_dim6,
				SV_dim7 => SV7_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s7
				);

	Kernel_rbf_8 : Kernel_rbf
	port map(	SV_dim0 => SV8_dim0,
				SV_dim1 => SV8_dim1,
				SV_dim2 => SV8_dim2,
				SV_dim3 => SV8_dim3,
				SV_dim4 => SV8_dim4,
				SV_dim5 => SV8_dim5,
				SV_dim6 => SV8_dim6,
				SV_dim7 => SV8_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s8
				);

	Kernel_rbf_9 : Kernel_rbf
	port map(	SV_dim0 => SV9_dim0,
				SV_dim1 => SV9_dim1,
				SV_dim2 => SV9_dim2,
				SV_dim3 => SV9_dim3,
				SV_dim4 => SV9_dim4,
				SV_dim5 => SV9_dim5,
				SV_dim6 => SV9_dim6,
				SV_dim7 => SV9_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s9
				);

	Kernel_rbf_10 : Kernel_rbf
	port map(	SV_dim0 => SV10_dim0,
				SV_dim1 => SV10_dim1,
				SV_dim2 => SV10_dim2,
				SV_dim3 => SV10_dim3,
				SV_dim4 => SV10_dim4,
				SV_dim5 => SV10_dim5,
				SV_dim6 => SV10_dim6,
				SV_dim7 => SV10_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s10
				);

	Kernel_rbf_11 : Kernel_rbf
	port map(	SV_dim0 => SV11_dim0,
				SV_dim1 => SV11_dim1,
				SV_dim2 => SV11_dim2,
				SV_dim3 => SV11_dim3,
				SV_dim4 => SV11_dim4,
				SV_dim5 => SV11_dim5,
				SV_dim6 => SV11_dim6,
				SV_dim7 => SV11_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s11
				);

	Kernel_rbf_12 : Kernel_rbf
	port map(	SV_dim0 => SV12_dim0,
				SV_dim1 => SV12_dim1,
				SV_dim2 => SV12_dim2,
				SV_dim3 => SV12_dim3,
				SV_dim4 => SV12_dim4,
				SV_dim5 => SV12_dim5,
				SV_dim6 => SV12_dim6,
				SV_dim7 => SV12_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s12
				);

	Kernel_rbf_13 : Kernel_rbf
	port map(	SV_dim0 => SV13_dim0,
				SV_dim1 => SV13_dim1,
				SV_dim2 => SV13_dim2,
				SV_dim3 => SV13_dim3,
				SV_dim4 => SV13_dim4,
				SV_dim5 => SV13_dim5,
				SV_dim6 => SV13_dim6,
				SV_dim7 => SV13_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s13
				);

	Kernel_rbf_14 : Kernel_rbf
	port map(	SV_dim0 => SV14_dim0,
				SV_dim1 => SV14_dim1,
				SV_dim2 => SV14_dim2,
				SV_dim3 => SV14_dim3,
				SV_dim4 => SV14_dim4,
				SV_dim5 => SV14_dim5,
				SV_dim6 => SV14_dim6,
				SV_dim7 => SV14_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s14
				);

	Kernel_rbf_15 : Kernel_rbf
	port map(	SV_dim0 => SV15_dim0,
				SV_dim1 => SV15_dim1,
				SV_dim2 => SV15_dim2,
				SV_dim3 => SV15_dim3,
				SV_dim4 => SV15_dim4,
				SV_dim5 => SV15_dim5,
				SV_dim6 => SV15_dim6,
				SV_dim7 => SV15_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s15
				);

	Kernel_rbf_16 : Kernel_rbf
	port map(	SV_dim0 => SV16_dim0,
				SV_dim1 => SV16_dim1,
				SV_dim2 => SV16_dim2,
				SV_dim3 => SV16_dim3,
				SV_dim4 => SV16_dim4,
				SV_dim5 => SV16_dim5,
				SV_dim6 => SV16_dim6,
				SV_dim7 => SV16_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s16
				);

	Kernel_rbf_17 : Kernel_rbf
	port map(	SV_dim0 => SV17_dim0,
				SV_dim1 => SV17_dim1,
				SV_dim2 => SV17_dim2,
				SV_dim3 => SV17_dim3,
				SV_dim4 => SV17_dim4,
				SV_dim5 => SV17_dim5,
				SV_dim6 => SV17_dim6,
				SV_dim7 => SV17_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s17
				);

	Kernel_rbf_18 : Kernel_rbf
	port map(	SV_dim0 => SV18_dim0,
				SV_dim1 => SV18_dim1,
				SV_dim2 => SV18_dim2,
				SV_dim3 => SV18_dim3,
				SV_dim4 => SV18_dim4,
				SV_dim5 => SV18_dim5,
				SV_dim6 => SV18_dim6,
				SV_dim7 => SV18_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s18
				);

	Kernel_rbf_19 : Kernel_rbf
	port map(	SV_dim0 => SV19_dim0,
				SV_dim1 => SV19_dim1,
				SV_dim2 => SV19_dim2,
				SV_dim3 => SV19_dim3,
				SV_dim4 => SV19_dim4,
				SV_dim5 => SV19_dim5,
				SV_dim6 => SV19_dim6,
				SV_dim7 => SV19_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s19
				);

	Kernel_rbf_20 : Kernel_rbf
	port map(	SV_dim0 => SV20_dim0,
				SV_dim1 => SV20_dim1,
				SV_dim2 => SV20_dim2,
				SV_dim3 => SV20_dim3,
				SV_dim4 => SV20_dim4,
				SV_dim5 => SV20_dim5,
				SV_dim6 => SV20_dim6,
				SV_dim7 => SV20_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s20
				);

	Kernel_rbf_21 : Kernel_rbf
	port map(	SV_dim0 => SV21_dim0,
				SV_dim1 => SV21_dim1,
				SV_dim2 => SV21_dim2,
				SV_dim3 => SV21_dim3,
				SV_dim4 => SV21_dim4,
				SV_dim5 => SV21_dim5,
				SV_dim6 => SV21_dim6,
				SV_dim7 => SV21_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s21
				);

	Kernel_rbf_22 : Kernel_rbf
	port map(	SV_dim0 => SV22_dim0,
				SV_dim1 => SV22_dim1,
				SV_dim2 => SV22_dim2,
				SV_dim3 => SV22_dim3,
				SV_dim4 => SV22_dim4,
				SV_dim5 => SV22_dim5,
				SV_dim6 => SV22_dim6,
				SV_dim7 => SV22_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s22
				);

	Kernel_rbf_23 : Kernel_rbf
	port map(	SV_dim0 => SV23_dim0,
				SV_dim1 => SV23_dim1,
				SV_dim2 => SV23_dim2,
				SV_dim3 => SV23_dim3,
				SV_dim4 => SV23_dim4,
				SV_dim5 => SV23_dim5,
				SV_dim6 => SV23_dim6,
				SV_dim7 => SV23_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s23
				);

	Kernel_rbf_24 : Kernel_rbf
	port map(	SV_dim0 => SV24_dim0,
				SV_dim1 => SV24_dim1,
				SV_dim2 => SV24_dim2,
				SV_dim3 => SV24_dim3,
				SV_dim4 => SV24_dim4,
				SV_dim5 => SV24_dim5,
				SV_dim6 => SV24_dim6,
				SV_dim7 => SV24_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s24
				);

	Kernel_rbf_25 : Kernel_rbf
	port map(	SV_dim0 => SV25_dim0,
				SV_dim1 => SV25_dim1,
				SV_dim2 => SV25_dim2,
				SV_dim3 => SV25_dim3,
				SV_dim4 => SV25_dim4,
				SV_dim5 => SV25_dim5,
				SV_dim6 => SV25_dim6,
				SV_dim7 => SV25_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s25
				);

	Kernel_rbf_26 : Kernel_rbf
	port map(	SV_dim0 => SV26_dim0,
				SV_dim1 => SV26_dim1,
				SV_dim2 => SV26_dim2,
				SV_dim3 => SV26_dim3,
				SV_dim4 => SV26_dim4,
				SV_dim5 => SV26_dim5,
				SV_dim6 => SV26_dim6,
				SV_dim7 => SV26_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s26
				);

	Kernel_rbf_27 : Kernel_rbf
	port map(	SV_dim0 => SV27_dim0,
				SV_dim1 => SV27_dim1,
				SV_dim2 => SV27_dim2,
				SV_dim3 => SV27_dim3,
				SV_dim4 => SV27_dim4,
				SV_dim5 => SV27_dim5,
				SV_dim6 => SV27_dim6,
				SV_dim7 => SV27_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s27
				);

	Kernel_rbf_28 : Kernel_rbf
	port map(	SV_dim0 => SV28_dim0,
				SV_dim1 => SV28_dim1,
				SV_dim2 => SV28_dim2,
				SV_dim3 => SV28_dim3,
				SV_dim4 => SV28_dim4,
				SV_dim5 => SV28_dim5,
				SV_dim6 => SV28_dim6,
				SV_dim7 => SV28_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s28
				);

	Kernel_rbf_29 : Kernel_rbf
	port map(	SV_dim0 => SV29_dim0,
				SV_dim1 => SV29_dim1,
				SV_dim2 => SV29_dim2,
				SV_dim3 => SV29_dim3,
				SV_dim4 => SV29_dim4,
				SV_dim5 => SV29_dim5,
				SV_dim6 => SV29_dim6,
				SV_dim7 => SV29_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s29
				);

	Kernel_rbf_30 : Kernel_rbf
	port map(	SV_dim0 => SV30_dim0,
				SV_dim1 => SV30_dim1,
				SV_dim2 => SV30_dim2,
				SV_dim3 => SV30_dim3,
				SV_dim4 => SV30_dim4,
				SV_dim5 => SV30_dim5,
				SV_dim6 => SV30_dim6,
				SV_dim7 => SV30_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s30
				);

	Kernel_rbf_31 : Kernel_rbf
	port map(	SV_dim0 => SV31_dim0,
				SV_dim1 => SV31_dim1,
				SV_dim2 => SV31_dim2,
				SV_dim3 => SV31_dim3,
				SV_dim4 => SV31_dim4,
				SV_dim5 => SV31_dim5,
				SV_dim6 => SV31_dim6,
				SV_dim7 => SV31_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s31
				);

	Kernel_rbf_32 : Kernel_rbf
	port map(	SV_dim0 => SV32_dim0,
				SV_dim1 => SV32_dim1,
				SV_dim2 => SV32_dim2,
				SV_dim3 => SV32_dim3,
				SV_dim4 => SV32_dim4,
				SV_dim5 => SV32_dim5,
				SV_dim6 => SV32_dim6,
				SV_dim7 => SV32_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s32
				);

	Kernel_rbf_33 : Kernel_rbf
	port map(	SV_dim0 => SV33_dim0,
				SV_dim1 => SV33_dim1,
				SV_dim2 => SV33_dim2,
				SV_dim3 => SV33_dim3,
				SV_dim4 => SV33_dim4,
				SV_dim5 => SV33_dim5,
				SV_dim6 => SV33_dim6,
				SV_dim7 => SV33_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s33
				);

	Kernel_rbf_34 : Kernel_rbf
	port map(	SV_dim0 => SV34_dim0,
				SV_dim1 => SV34_dim1,
				SV_dim2 => SV34_dim2,
				SV_dim3 => SV34_dim3,
				SV_dim4 => SV34_dim4,
				SV_dim5 => SV34_dim5,
				SV_dim6 => SV34_dim6,
				SV_dim7 => SV34_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s34
				);

	Kernel_rbf_35 : Kernel_rbf
	port map(	SV_dim0 => SV35_dim0,
				SV_dim1 => SV35_dim1,
				SV_dim2 => SV35_dim2,
				SV_dim3 => SV35_dim3,
				SV_dim4 => SV35_dim4,
				SV_dim5 => SV35_dim5,
				SV_dim6 => SV35_dim6,
				SV_dim7 => SV35_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s35
				);

	Kernel_rbf_36 : Kernel_rbf
	port map(	SV_dim0 => SV36_dim0,
				SV_dim1 => SV36_dim1,
				SV_dim2 => SV36_dim2,
				SV_dim3 => SV36_dim3,
				SV_dim4 => SV36_dim4,
				SV_dim5 => SV36_dim5,
				SV_dim6 => SV36_dim6,
				SV_dim7 => SV36_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s36
				);

	Kernel_rbf_37 : Kernel_rbf
	port map(	SV_dim0 => SV37_dim0,
				SV_dim1 => SV37_dim1,
				SV_dim2 => SV37_dim2,
				SV_dim3 => SV37_dim3,
				SV_dim4 => SV37_dim4,
				SV_dim5 => SV37_dim5,
				SV_dim6 => SV37_dim6,
				SV_dim7 => SV37_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s37
				);

	Kernel_rbf_38 : Kernel_rbf
	port map(	SV_dim0 => SV38_dim0,
				SV_dim1 => SV38_dim1,
				SV_dim2 => SV38_dim2,
				SV_dim3 => SV38_dim3,
				SV_dim4 => SV38_dim4,
				SV_dim5 => SV38_dim5,
				SV_dim6 => SV38_dim6,
				SV_dim7 => SV38_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s38
				);

	Kernel_rbf_39 : Kernel_rbf
	port map(	SV_dim0 => SV39_dim0,
				SV_dim1 => SV39_dim1,
				SV_dim2 => SV39_dim2,
				SV_dim3 => SV39_dim3,
				SV_dim4 => SV39_dim4,
				SV_dim5 => SV39_dim5,
				SV_dim6 => SV39_dim6,
				SV_dim7 => SV39_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s39
				);

	Kernel_rbf_40 : Kernel_rbf
	port map(	SV_dim0 => SV40_dim0,
				SV_dim1 => SV40_dim1,
				SV_dim2 => SV40_dim2,
				SV_dim3 => SV40_dim3,
				SV_dim4 => SV40_dim4,
				SV_dim5 => SV40_dim5,
				SV_dim6 => SV40_dim6,
				SV_dim7 => SV40_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s40
				);

	Kernel_rbf_41 : Kernel_rbf
	port map(	SV_dim0 => SV41_dim0,
				SV_dim1 => SV41_dim1,
				SV_dim2 => SV41_dim2,
				SV_dim3 => SV41_dim3,
				SV_dim4 => SV41_dim4,
				SV_dim5 => SV41_dim5,
				SV_dim6 => SV41_dim6,
				SV_dim7 => SV41_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s41
				);

	Kernel_rbf_42 : Kernel_rbf
	port map(	SV_dim0 => SV42_dim0,
				SV_dim1 => SV42_dim1,
				SV_dim2 => SV42_dim2,
				SV_dim3 => SV42_dim3,
				SV_dim4 => SV42_dim4,
				SV_dim5 => SV42_dim5,
				SV_dim6 => SV42_dim6,
				SV_dim7 => SV42_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s42
				);

	Kernel_rbf_43 : Kernel_rbf
	port map(	SV_dim0 => SV43_dim0,
				SV_dim1 => SV43_dim1,
				SV_dim2 => SV43_dim2,
				SV_dim3 => SV43_dim3,
				SV_dim4 => SV43_dim4,
				SV_dim5 => SV43_dim5,
				SV_dim6 => SV43_dim6,
				SV_dim7 => SV43_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s43
				);

	Kernel_rbf_44 : Kernel_rbf
	port map(	SV_dim0 => SV44_dim0,
				SV_dim1 => SV44_dim1,
				SV_dim2 => SV44_dim2,
				SV_dim3 => SV44_dim3,
				SV_dim4 => SV44_dim4,
				SV_dim5 => SV44_dim5,
				SV_dim6 => SV44_dim6,
				SV_dim7 => SV44_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s44
				);

	Kernel_rbf_45 : Kernel_rbf
	port map(	SV_dim0 => SV45_dim0,
				SV_dim1 => SV45_dim1,
				SV_dim2 => SV45_dim2,
				SV_dim3 => SV45_dim3,
				SV_dim4 => SV45_dim4,
				SV_dim5 => SV45_dim5,
				SV_dim6 => SV45_dim6,
				SV_dim7 => SV45_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s45
				);

	Kernel_rbf_46 : Kernel_rbf
	port map(	SV_dim0 => SV46_dim0,
				SV_dim1 => SV46_dim1,
				SV_dim2 => SV46_dim2,
				SV_dim3 => SV46_dim3,
				SV_dim4 => SV46_dim4,
				SV_dim5 => SV46_dim5,
				SV_dim6 => SV46_dim6,
				SV_dim7 => SV46_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s46
				);

	Kernel_rbf_47 : Kernel_rbf
	port map(	SV_dim0 => SV47_dim0,
				SV_dim1 => SV47_dim1,
				SV_dim2 => SV47_dim2,
				SV_dim3 => SV47_dim3,
				SV_dim4 => SV47_dim4,
				SV_dim5 => SV47_dim5,
				SV_dim6 => SV47_dim6,
				SV_dim7 => SV47_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s47
				);

	Kernel_rbf_48 : Kernel_rbf
	port map(	SV_dim0 => SV48_dim0,
				SV_dim1 => SV48_dim1,
				SV_dim2 => SV48_dim2,
				SV_dim3 => SV48_dim3,
				SV_dim4 => SV48_dim4,
				SV_dim5 => SV48_dim5,
				SV_dim6 => SV48_dim6,
				SV_dim7 => SV48_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s48
				);

	Kernel_rbf_49 : Kernel_rbf
	port map(	SV_dim0 => SV49_dim0,
				SV_dim1 => SV49_dim1,
				SV_dim2 => SV49_dim2,
				SV_dim3 => SV49_dim3,
				SV_dim4 => SV49_dim4,
				SV_dim5 => SV49_dim5,
				SV_dim6 => SV49_dim6,
				SV_dim7 => SV49_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s49
				);

	Kernel_rbf_50 : Kernel_rbf
	port map(	SV_dim0 => SV50_dim0,
				SV_dim1 => SV50_dim1,
				SV_dim2 => SV50_dim2,
				SV_dim3 => SV50_dim3,
				SV_dim4 => SV50_dim4,
				SV_dim5 => SV50_dim5,
				SV_dim6 => SV50_dim6,
				SV_dim7 => SV50_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s50
				);

	Kernel_rbf_51 : Kernel_rbf
	port map(	SV_dim0 => SV51_dim0,
				SV_dim1 => SV51_dim1,
				SV_dim2 => SV51_dim2,
				SV_dim3 => SV51_dim3,
				SV_dim4 => SV51_dim4,
				SV_dim5 => SV51_dim5,
				SV_dim6 => SV51_dim6,
				SV_dim7 => SV51_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s51
				);

	Kernel_rbf_52 : Kernel_rbf
	port map(	SV_dim0 => SV52_dim0,
				SV_dim1 => SV52_dim1,
				SV_dim2 => SV52_dim2,
				SV_dim3 => SV52_dim3,
				SV_dim4 => SV52_dim4,
				SV_dim5 => SV52_dim5,
				SV_dim6 => SV52_dim6,
				SV_dim7 => SV52_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s52
				);

	Kernel_rbf_53 : Kernel_rbf
	port map(	SV_dim0 => SV53_dim0,
				SV_dim1 => SV53_dim1,
				SV_dim2 => SV53_dim2,
				SV_dim3 => SV53_dim3,
				SV_dim4 => SV53_dim4,
				SV_dim5 => SV53_dim5,
				SV_dim6 => SV53_dim6,
				SV_dim7 => SV53_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s53
				);

	Kernel_rbf_54 : Kernel_rbf
	port map(	SV_dim0 => SV54_dim0,
				SV_dim1 => SV54_dim1,
				SV_dim2 => SV54_dim2,
				SV_dim3 => SV54_dim3,
				SV_dim4 => SV54_dim4,
				SV_dim5 => SV54_dim5,
				SV_dim6 => SV54_dim6,
				SV_dim7 => SV54_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s54
				);

	Kernel_rbf_55 : Kernel_rbf
	port map(	SV_dim0 => SV55_dim0,
				SV_dim1 => SV55_dim1,
				SV_dim2 => SV55_dim2,
				SV_dim3 => SV55_dim3,
				SV_dim4 => SV55_dim4,
				SV_dim5 => SV55_dim5,
				SV_dim6 => SV55_dim6,
				SV_dim7 => SV55_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s55
				);

	Kernel_rbf_56 : Kernel_rbf
	port map(	SV_dim0 => SV56_dim0,
				SV_dim1 => SV56_dim1,
				SV_dim2 => SV56_dim2,
				SV_dim3 => SV56_dim3,
				SV_dim4 => SV56_dim4,
				SV_dim5 => SV56_dim5,
				SV_dim6 => SV56_dim6,
				SV_dim7 => SV56_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s56
				);

	Kernel_rbf_57 : Kernel_rbf
	port map(	SV_dim0 => SV57_dim0,
				SV_dim1 => SV57_dim1,
				SV_dim2 => SV57_dim2,
				SV_dim3 => SV57_dim3,
				SV_dim4 => SV57_dim4,
				SV_dim5 => SV57_dim5,
				SV_dim6 => SV57_dim6,
				SV_dim7 => SV57_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s57
				);

	Kernel_rbf_58 : Kernel_rbf
	port map(	SV_dim0 => SV58_dim0,
				SV_dim1 => SV58_dim1,
				SV_dim2 => SV58_dim2,
				SV_dim3 => SV58_dim3,
				SV_dim4 => SV58_dim4,
				SV_dim5 => SV58_dim5,
				SV_dim6 => SV58_dim6,
				SV_dim7 => SV58_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s58
				);

	Kernel_rbf_59 : Kernel_rbf
	port map(	SV_dim0 => SV59_dim0,
				SV_dim1 => SV59_dim1,
				SV_dim2 => SV59_dim2,
				SV_dim3 => SV59_dim3,
				SV_dim4 => SV59_dim4,
				SV_dim5 => SV59_dim5,
				SV_dim6 => SV59_dim6,
				SV_dim7 => SV59_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s59
				);

	Kernel_rbf_60 : Kernel_rbf
	port map(	SV_dim0 => SV60_dim0,
				SV_dim1 => SV60_dim1,
				SV_dim2 => SV60_dim2,
				SV_dim3 => SV60_dim3,
				SV_dim4 => SV60_dim4,
				SV_dim5 => SV60_dim5,
				SV_dim6 => SV60_dim6,
				SV_dim7 => SV60_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s60
				);

	Kernel_rbf_61 : Kernel_rbf
	port map(	SV_dim0 => SV61_dim0,
				SV_dim1 => SV61_dim1,
				SV_dim2 => SV61_dim2,
				SV_dim3 => SV61_dim3,
				SV_dim4 => SV61_dim4,
				SV_dim5 => SV61_dim5,
				SV_dim6 => SV61_dim6,
				SV_dim7 => SV61_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s61
				);

	Kernel_rbf_62 : Kernel_rbf
	port map(	SV_dim0 => SV62_dim0,
				SV_dim1 => SV62_dim1,
				SV_dim2 => SV62_dim2,
				SV_dim3 => SV62_dim3,
				SV_dim4 => SV62_dim4,
				SV_dim5 => SV62_dim5,
				SV_dim6 => SV62_dim6,
				SV_dim7 => SV62_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s62
				);

	Kernel_rbf_63 : Kernel_rbf
	port map(	SV_dim0 => SV63_dim0,
				SV_dim1 => SV63_dim1,
				SV_dim2 => SV63_dim2,
				SV_dim3 => SV63_dim3,
				SV_dim4 => SV63_dim4,
				SV_dim5 => SV63_dim5,
				SV_dim6 => SV63_dim6,
				SV_dim7 => SV63_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s63
				);

	Kernel_rbf_64 : Kernel_rbf
	port map(	SV_dim0 => SV64_dim0,
				SV_dim1 => SV64_dim1,
				SV_dim2 => SV64_dim2,
				SV_dim3 => SV64_dim3,
				SV_dim4 => SV64_dim4,
				SV_dim5 => SV64_dim5,
				SV_dim6 => SV64_dim6,
				SV_dim7 => SV64_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s64
				);

	Kernel_rbf_65 : Kernel_rbf
	port map(	SV_dim0 => SV65_dim0,
				SV_dim1 => SV65_dim1,
				SV_dim2 => SV65_dim2,
				SV_dim3 => SV65_dim3,
				SV_dim4 => SV65_dim4,
				SV_dim5 => SV65_dim5,
				SV_dim6 => SV65_dim6,
				SV_dim7 => SV65_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s65
				);

	Kernel_rbf_66 : Kernel_rbf
	port map(	SV_dim0 => SV66_dim0,
				SV_dim1 => SV66_dim1,
				SV_dim2 => SV66_dim2,
				SV_dim3 => SV66_dim3,
				SV_dim4 => SV66_dim4,
				SV_dim5 => SV66_dim5,
				SV_dim6 => SV66_dim6,
				SV_dim7 => SV66_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s66
				);

	Kernel_rbf_67 : Kernel_rbf
	port map(	SV_dim0 => SV67_dim0,
				SV_dim1 => SV67_dim1,
				SV_dim2 => SV67_dim2,
				SV_dim3 => SV67_dim3,
				SV_dim4 => SV67_dim4,
				SV_dim5 => SV67_dim5,
				SV_dim6 => SV67_dim6,
				SV_dim7 => SV67_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s67
				);

	Kernel_rbf_68 : Kernel_rbf
	port map(	SV_dim0 => SV68_dim0,
				SV_dim1 => SV68_dim1,
				SV_dim2 => SV68_dim2,
				SV_dim3 => SV68_dim3,
				SV_dim4 => SV68_dim4,
				SV_dim5 => SV68_dim5,
				SV_dim6 => SV68_dim6,
				SV_dim7 => SV68_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s68
				);

	Kernel_rbf_69 : Kernel_rbf
	port map(	SV_dim0 => SV69_dim0,
				SV_dim1 => SV69_dim1,
				SV_dim2 => SV69_dim2,
				SV_dim3 => SV69_dim3,
				SV_dim4 => SV69_dim4,
				SV_dim5 => SV69_dim5,
				SV_dim6 => SV69_dim6,
				SV_dim7 => SV69_dim7,
				test_data_dim0 => test_data_dim00,
				test_data_dim1 => test_data_dim01,
				test_data_dim2 => test_data_dim02,
				test_data_dim3 => test_data_dim03,
				test_data_dim4 => test_data_dim04,
				test_data_dim5 => test_data_dim05,
				test_data_dim6 => test_data_dim06,
				test_data_dim7 => test_data_dim07,
				gamma => gamma,
				output => Kernel_rbf_output_s69
				);

	Multiplier_Signed_12bits_0 : Multiplier_Signed_12bits
	port map(	input_a => SV0_alphaY,
				input_b => '0' & Kernel_rbf_output_s0,
				output => multi_s0
				);

	Multiplier_Signed_12bits_1 : Multiplier_Signed_12bits
	port map(	input_a => SV1_alphaY,
				input_b => '0' & Kernel_rbf_output_s1,
				output => multi_s1
				);

	Multiplier_Signed_12bits_2 : Multiplier_Signed_12bits
	port map(	input_a => SV2_alphaY,
				input_b => '0' & Kernel_rbf_output_s2,
				output => multi_s2
				);

	Multiplier_Signed_12bits_3 : Multiplier_Signed_12bits
	port map(	input_a => SV3_alphaY,
				input_b => '0' & Kernel_rbf_output_s3,
				output => multi_s3
				);

	Multiplier_Signed_12bits_4 : Multiplier_Signed_12bits
	port map(	input_a => SV4_alphaY,
				input_b => '0' & Kernel_rbf_output_s4,
				output => multi_s4
				);

	Multiplier_Signed_12bits_5 : Multiplier_Signed_12bits
	port map(	input_a => SV5_alphaY,
				input_b => '0' & Kernel_rbf_output_s5,
				output => multi_s5
				);

	Multiplier_Signed_12bits_6 : Multiplier_Signed_12bits
	port map(	input_a => SV6_alphaY,
				input_b => '0' & Kernel_rbf_output_s6,
				output => multi_s6
				);

	Multiplier_Signed_12bits_7 : Multiplier_Signed_12bits
	port map(	input_a => SV7_alphaY,
				input_b => '0' & Kernel_rbf_output_s7,
				output => multi_s7
				);

	Multiplier_Signed_12bits_8 : Multiplier_Signed_12bits
	port map(	input_a => SV8_alphaY,
				input_b => '0' & Kernel_rbf_output_s8,
				output => multi_s8
				);

	Multiplier_Signed_12bits_9 : Multiplier_Signed_12bits
	port map(	input_a => SV9_alphaY,
				input_b => '0' & Kernel_rbf_output_s9,
				output => multi_s9
				);

	Multiplier_Signed_12bits_10 : Multiplier_Signed_12bits
	port map(	input_a => SV10_alphaY,
				input_b => '0' & Kernel_rbf_output_s10,
				output => multi_s10
				);

	Multiplier_Signed_12bits_11 : Multiplier_Signed_12bits
	port map(	input_a => SV11_alphaY,
				input_b => '0' & Kernel_rbf_output_s11,
				output => multi_s11
				);

	Multiplier_Signed_12bits_12 : Multiplier_Signed_12bits
	port map(	input_a => SV12_alphaY,
				input_b => '0' & Kernel_rbf_output_s12,
				output => multi_s12
				);

	Multiplier_Signed_12bits_13 : Multiplier_Signed_12bits
	port map(	input_a => SV13_alphaY,
				input_b => '0' & Kernel_rbf_output_s13,
				output => multi_s13
				);

	Multiplier_Signed_12bits_14 : Multiplier_Signed_12bits
	port map(	input_a => SV14_alphaY,
				input_b => '0' & Kernel_rbf_output_s14,
				output => multi_s14
				);

	Multiplier_Signed_12bits_15 : Multiplier_Signed_12bits
	port map(	input_a => SV15_alphaY,
				input_b => '0' & Kernel_rbf_output_s15,
				output => multi_s15
				);

	Multiplier_Signed_12bits_16 : Multiplier_Signed_12bits
	port map(	input_a => SV16_alphaY,
				input_b => '0' & Kernel_rbf_output_s16,
				output => multi_s16
				);

	Multiplier_Signed_12bits_17 : Multiplier_Signed_12bits
	port map(	input_a => SV17_alphaY,
				input_b => '0' & Kernel_rbf_output_s17,
				output => multi_s17
				);

	Multiplier_Signed_12bits_18 : Multiplier_Signed_12bits
	port map(	input_a => SV18_alphaY,
				input_b => '0' & Kernel_rbf_output_s18,
				output => multi_s18
				);

	Multiplier_Signed_12bits_19 : Multiplier_Signed_12bits
	port map(	input_a => SV19_alphaY,
				input_b => '0' & Kernel_rbf_output_s19,
				output => multi_s19
				);

	Multiplier_Signed_12bits_20 : Multiplier_Signed_12bits
	port map(	input_a => SV20_alphaY,
				input_b => '0' & Kernel_rbf_output_s20,
				output => multi_s20
				);

	Multiplier_Signed_12bits_21 : Multiplier_Signed_12bits
	port map(	input_a => SV21_alphaY,
				input_b => '0' & Kernel_rbf_output_s21,
				output => multi_s21
				);

	Multiplier_Signed_12bits_22 : Multiplier_Signed_12bits
	port map(	input_a => SV22_alphaY,
				input_b => '0' & Kernel_rbf_output_s22,
				output => multi_s22
				);

	Multiplier_Signed_12bits_23 : Multiplier_Signed_12bits
	port map(	input_a => SV23_alphaY,
				input_b => '0' & Kernel_rbf_output_s23,
				output => multi_s23
				);

	Multiplier_Signed_12bits_24 : Multiplier_Signed_12bits
	port map(	input_a => SV24_alphaY,
				input_b => '0' & Kernel_rbf_output_s24,
				output => multi_s24
				);

	Multiplier_Signed_12bits_25 : Multiplier_Signed_12bits
	port map(	input_a => SV25_alphaY,
				input_b => '0' & Kernel_rbf_output_s25,
				output => multi_s25
				);

	Multiplier_Signed_12bits_26 : Multiplier_Signed_12bits
	port map(	input_a => SV26_alphaY,
				input_b => '0' & Kernel_rbf_output_s26,
				output => multi_s26
				);

	Multiplier_Signed_12bits_27 : Multiplier_Signed_12bits
	port map(	input_a => SV27_alphaY,
				input_b => '0' & Kernel_rbf_output_s27,
				output => multi_s27
				);

	Multiplier_Signed_12bits_28 : Multiplier_Signed_12bits
	port map(	input_a => SV28_alphaY,
				input_b => '0' & Kernel_rbf_output_s28,
				output => multi_s28
				);

	Multiplier_Signed_12bits_29 : Multiplier_Signed_12bits
	port map(	input_a => SV29_alphaY,
				input_b => '0' & Kernel_rbf_output_s29,
				output => multi_s29
				);

	Multiplier_Signed_12bits_30 : Multiplier_Signed_12bits
	port map(	input_a => SV30_alphaY,
				input_b => '0' & Kernel_rbf_output_s30,
				output => multi_s30
				);

	Multiplier_Signed_12bits_31 : Multiplier_Signed_12bits
	port map(	input_a => SV31_alphaY,
				input_b => '0' & Kernel_rbf_output_s31,
				output => multi_s31
				);

	Multiplier_Signed_12bits_32 : Multiplier_Signed_12bits
	port map(	input_a => SV32_alphaY,
				input_b => '0' & Kernel_rbf_output_s32,
				output => multi_s32
				);

	Multiplier_Signed_12bits_33 : Multiplier_Signed_12bits
	port map(	input_a => SV33_alphaY,
				input_b => '0' & Kernel_rbf_output_s33,
				output => multi_s33
				);

	Multiplier_Signed_12bits_34 : Multiplier_Signed_12bits
	port map(	input_a => SV34_alphaY,
				input_b => '0' & Kernel_rbf_output_s34,
				output => multi_s34
				);

	Multiplier_Signed_12bits_35 : Multiplier_Signed_12bits
	port map(	input_a => SV35_alphaY,
				input_b => '0' & Kernel_rbf_output_s35,
				output => multi_s35
				);

	Multiplier_Signed_12bits_36 : Multiplier_Signed_12bits
	port map(	input_a => SV36_alphaY,
				input_b => '0' & Kernel_rbf_output_s36,
				output => multi_s36
				);

	Multiplier_Signed_12bits_37 : Multiplier_Signed_12bits
	port map(	input_a => SV37_alphaY,
				input_b => '0' & Kernel_rbf_output_s37,
				output => multi_s37
				);

	Multiplier_Signed_12bits_38 : Multiplier_Signed_12bits
	port map(	input_a => SV38_alphaY,
				input_b => '0' & Kernel_rbf_output_s38,
				output => multi_s38
				);

	Multiplier_Signed_12bits_39 : Multiplier_Signed_12bits
	port map(	input_a => SV39_alphaY,
				input_b => '0' & Kernel_rbf_output_s39,
				output => multi_s39
				);

	Multiplier_Signed_12bits_40 : Multiplier_Signed_12bits
	port map(	input_a => SV40_alphaY,
				input_b => '0' & Kernel_rbf_output_s40,
				output => multi_s40
				);

	Multiplier_Signed_12bits_41 : Multiplier_Signed_12bits
	port map(	input_a => SV41_alphaY,
				input_b => '0' & Kernel_rbf_output_s41,
				output => multi_s41
				);

	Multiplier_Signed_12bits_42 : Multiplier_Signed_12bits
	port map(	input_a => SV42_alphaY,
				input_b => '0' & Kernel_rbf_output_s42,
				output => multi_s42
				);

	Multiplier_Signed_12bits_43 : Multiplier_Signed_12bits
	port map(	input_a => SV43_alphaY,
				input_b => '0' & Kernel_rbf_output_s43,
				output => multi_s43
				);

	Multiplier_Signed_12bits_44 : Multiplier_Signed_12bits
	port map(	input_a => SV44_alphaY,
				input_b => '0' & Kernel_rbf_output_s44,
				output => multi_s44
				);

	Multiplier_Signed_12bits_45 : Multiplier_Signed_12bits
	port map(	input_a => SV45_alphaY,
				input_b => '0' & Kernel_rbf_output_s45,
				output => multi_s45
				);

	Multiplier_Signed_12bits_46 : Multiplier_Signed_12bits
	port map(	input_a => SV46_alphaY,
				input_b => '0' & Kernel_rbf_output_s46,
				output => multi_s46
				);

	Multiplier_Signed_12bits_47 : Multiplier_Signed_12bits
	port map(	input_a => SV47_alphaY,
				input_b => '0' & Kernel_rbf_output_s47,
				output => multi_s47
				);

	Multiplier_Signed_12bits_48 : Multiplier_Signed_12bits
	port map(	input_a => SV48_alphaY,
				input_b => '0' & Kernel_rbf_output_s48,
				output => multi_s48
				);

	Multiplier_Signed_12bits_49 : Multiplier_Signed_12bits
	port map(	input_a => SV49_alphaY,
				input_b => '0' & Kernel_rbf_output_s49,
				output => multi_s49
				);

	Multiplier_Signed_12bits_50 : Multiplier_Signed_12bits
	port map(	input_a => SV50_alphaY,
				input_b => '0' & Kernel_rbf_output_s50,
				output => multi_s50
				);

	Multiplier_Signed_12bits_51 : Multiplier_Signed_12bits
	port map(	input_a => SV51_alphaY,
				input_b => '0' & Kernel_rbf_output_s51,
				output => multi_s51
				);

	Multiplier_Signed_12bits_52 : Multiplier_Signed_12bits
	port map(	input_a => SV52_alphaY,
				input_b => '0' & Kernel_rbf_output_s52,
				output => multi_s52
				);

	Multiplier_Signed_12bits_53 : Multiplier_Signed_12bits
	port map(	input_a => SV53_alphaY,
				input_b => '0' & Kernel_rbf_output_s53,
				output => multi_s53
				);

	Multiplier_Signed_12bits_54 : Multiplier_Signed_12bits
	port map(	input_a => SV54_alphaY,
				input_b => '0' & Kernel_rbf_output_s54,
				output => multi_s54
				);

	Multiplier_Signed_12bits_55 : Multiplier_Signed_12bits
	port map(	input_a => SV55_alphaY,
				input_b => '0' & Kernel_rbf_output_s55,
				output => multi_s55
				);

	Multiplier_Signed_12bits_56 : Multiplier_Signed_12bits
	port map(	input_a => SV56_alphaY,
				input_b => '0' & Kernel_rbf_output_s56,
				output => multi_s56
				);

	Multiplier_Signed_12bits_57 : Multiplier_Signed_12bits
	port map(	input_a => SV57_alphaY,
				input_b => '0' & Kernel_rbf_output_s57,
				output => multi_s57
				);

	Multiplier_Signed_12bits_58 : Multiplier_Signed_12bits
	port map(	input_a => SV58_alphaY,
				input_b => '0' & Kernel_rbf_output_s58,
				output => multi_s58
				);

	Multiplier_Signed_12bits_59 : Multiplier_Signed_12bits
	port map(	input_a => SV59_alphaY,
				input_b => '0' & Kernel_rbf_output_s59,
				output => multi_s59
				);

	Multiplier_Signed_12bits_60 : Multiplier_Signed_12bits
	port map(	input_a => SV60_alphaY,
				input_b => '0' & Kernel_rbf_output_s60,
				output => multi_s60
				);

	Multiplier_Signed_12bits_61 : Multiplier_Signed_12bits
	port map(	input_a => SV61_alphaY,
				input_b => '0' & Kernel_rbf_output_s61,
				output => multi_s61
				);

	Multiplier_Signed_12bits_62 : Multiplier_Signed_12bits
	port map(	input_a => SV62_alphaY,
				input_b => '0' & Kernel_rbf_output_s62,
				output => multi_s62
				);

	Multiplier_Signed_12bits_63 : Multiplier_Signed_12bits
	port map(	input_a => SV63_alphaY,
				input_b => '0' & Kernel_rbf_output_s63,
				output => multi_s63
				);

	Multiplier_Signed_12bits_64 : Multiplier_Signed_12bits
	port map(	input_a => SV64_alphaY,
				input_b => '0' & Kernel_rbf_output_s64,
				output => multi_s64
				);

	Multiplier_Signed_12bits_65 : Multiplier_Signed_12bits
	port map(	input_a => SV65_alphaY,
				input_b => '0' & Kernel_rbf_output_s65,
				output => multi_s65
				);

	Multiplier_Signed_12bits_66 : Multiplier_Signed_12bits
	port map(	input_a => SV66_alphaY,
				input_b => '0' & Kernel_rbf_output_s66,
				output => multi_s66
				);

	Multiplier_Signed_12bits_67 : Multiplier_Signed_12bits
	port map(	input_a => SV67_alphaY,
				input_b => '0' & Kernel_rbf_output_s67,
				output => multi_s67
				);

	Multiplier_Signed_12bits_68 : Multiplier_Signed_12bits
	port map(	input_a => SV68_alphaY,
				input_b => '0' & Kernel_rbf_output_s68,
				output => multi_s68
				);

	Multiplier_Signed_12bits_69 : Multiplier_Signed_12bits
	port map(	input_a => SV69_alphaY,
				input_b => '0' & Kernel_rbf_output_s69,
				output => multi_s69
				);

	Multiplier_Signed_12bits_70 : Multiplier_Signed_12bits
	port map(	input_a => SV70_alphaY,
				input_b => '0' & Kernel_rbf_output_s70,
				output => multi_s70
				);

	Adder_Signed_20bits_00 : Adder_Signed_20bits
	port map(	input_a => multi_s0,
				input_b => multi_s1,
				output => add_output_s00,
				overflow => add_overflow_s00
				);

	Adder_Signed_20bits_01 : Adder_Signed_20bits
	port map(	input_a => multi_s2,
				input_b => multi_s3,
				output => add_output_s01,
				overflow => add_overflow_s01
				);

	Adder_Signed_20bits_02 : Adder_Signed_20bits
	port map(	input_a => multi_s4,
				input_b => multi_s5,
				output => add_output_s02,
				overflow => add_overflow_s02
				);

	Adder_Signed_20bits_03 : Adder_Signed_20bits
	port map(	input_a => multi_s6,
				input_b => multi_s7,
				output => add_output_s03,
				overflow => add_overflow_s03
				);

	Adder_Signed_20bits_04 : Adder_Signed_20bits
	port map(	input_a => multi_s8,
				input_b => multi_s9,
				output => add_output_s04,
				overflow => add_overflow_s04
				);

	Adder_Signed_20bits_05 : Adder_Signed_20bits
	port map(	input_a => multi_s10,
				input_b => multi_s11,
				output => add_output_s05,
				overflow => add_overflow_s05
				);

	Adder_Signed_20bits_06 : Adder_Signed_20bits
	port map(	input_a => multi_s12,
				input_b => multi_s13,
				output => add_output_s06,
				overflow => add_overflow_s06
				);

	Adder_Signed_20bits_07 : Adder_Signed_20bits
	port map(	input_a => multi_s14,
				input_b => multi_s15,
				output => add_output_s07,
				overflow => add_overflow_s07
				);

	Adder_Signed_20bits_08 : Adder_Signed_20bits
	port map(	input_a => multi_s16,
				input_b => multi_s17,
				output => add_output_s08,
				overflow => add_overflow_s08
				);

	Adder_Signed_20bits_09 : Adder_Signed_20bits
	port map(	input_a => multi_s18,
				input_b => multi_s19,
				output => add_output_s09,
				overflow => add_overflow_s09
				);

	Adder_Signed_20bits_010 : Adder_Signed_20bits
	port map(	input_a => multi_s20,
				input_b => multi_s21,
				output => add_output_s010,
				overflow => add_overflow_s010
				);

	Adder_Signed_20bits_011 : Adder_Signed_20bits
	port map(	input_a => multi_s22,
				input_b => multi_s23,
				output => add_output_s011,
				overflow => add_overflow_s011
				);

	Adder_Signed_20bits_012 : Adder_Signed_20bits
	port map(	input_a => multi_s24,
				input_b => multi_s25,
				output => add_output_s012,
				overflow => add_overflow_s012
				);

	Adder_Signed_20bits_013 : Adder_Signed_20bits
	port map(	input_a => multi_s26,
				input_b => multi_s27,
				output => add_output_s013,
				overflow => add_overflow_s013
				);

	Adder_Signed_20bits_014 : Adder_Signed_20bits
	port map(	input_a => multi_s28,
				input_b => multi_s29,
				output => add_output_s014,
				overflow => add_overflow_s014
				);

	Adder_Signed_20bits_015 : Adder_Signed_20bits
	port map(	input_a => multi_s30,
				input_b => multi_s31,
				output => add_output_s015,
				overflow => add_overflow_s015
				);

	Adder_Signed_20bits_016 : Adder_Signed_20bits
	port map(	input_a => multi_s32,
				input_b => multi_s33,
				output => add_output_s016,
				overflow => add_overflow_s016
				);

	Adder_Signed_20bits_017 : Adder_Signed_20bits
	port map(	input_a => multi_s34,
				input_b => multi_s35,
				output => add_output_s017,
				overflow => add_overflow_s017
				);

	Adder_Signed_20bits_018 : Adder_Signed_20bits
	port map(	input_a => multi_s36,
				input_b => multi_s37,
				output => add_output_s018,
				overflow => add_overflow_s018
				);

	Adder_Signed_20bits_019 : Adder_Signed_20bits
	port map(	input_a => multi_s38,
				input_b => multi_s39,
				output => add_output_s019,
				overflow => add_overflow_s019
				);

	Adder_Signed_20bits_020 : Adder_Signed_20bits
	port map(	input_a => multi_s40,
				input_b => multi_s41,
				output => add_output_s020,
				overflow => add_overflow_s020
				);

	Adder_Signed_20bits_021 : Adder_Signed_20bits
	port map(	input_a => multi_s42,
				input_b => multi_s43,
				output => add_output_s021,
				overflow => add_overflow_s021
				);

	Adder_Signed_20bits_022 : Adder_Signed_20bits
	port map(	input_a => multi_s44,
				input_b => multi_s45,
				output => add_output_s022,
				overflow => add_overflow_s022
				);

	Adder_Signed_20bits_023 : Adder_Signed_20bits
	port map(	input_a => multi_s46,
				input_b => multi_s47,
				output => add_output_s023,
				overflow => add_overflow_s023
				);

	Adder_Signed_20bits_024 : Adder_Signed_20bits
	port map(	input_a => multi_s48,
				input_b => multi_s49,
				output => add_output_s024,
				overflow => add_overflow_s024
				);

	Adder_Signed_20bits_025 : Adder_Signed_20bits
	port map(	input_a => multi_s50,
				input_b => multi_s51,
				output => add_output_s025,
				overflow => add_overflow_s025
				);

	Adder_Signed_20bits_026 : Adder_Signed_20bits
	port map(	input_a => multi_s52,
				input_b => multi_s53,
				output => add_output_s026,
				overflow => add_overflow_s026
				);

	Adder_Signed_20bits_027 : Adder_Signed_20bits
	port map(	input_a => multi_s54,
				input_b => multi_s55,
				output => add_output_s027,
				overflow => add_overflow_s027
				);

	Adder_Signed_20bits_028 : Adder_Signed_20bits
	port map(	input_a => multi_s56,
				input_b => multi_s57,
				output => add_output_s028,
				overflow => add_overflow_s028
				);

	Adder_Signed_20bits_029 : Adder_Signed_20bits
	port map(	input_a => multi_s58,
				input_b => multi_s59,
				output => add_output_s029,
				overflow => add_overflow_s029
				);

	Adder_Signed_20bits_030 : Adder_Signed_20bits
	port map(	input_a => multi_s60,
				input_b => multi_s61,
				output => add_output_s030,
				overflow => add_overflow_s030
				);

	Adder_Signed_20bits_031 : Adder_Signed_20bits
	port map(	input_a => multi_s62,
				input_b => multi_s63,
				output => add_output_s031,
				overflow => add_overflow_s031
				);

	Adder_Signed_20bits_032 : Adder_Signed_20bits
	port map(	input_a => multi_s64,
				input_b => multi_s65,
				output => add_output_s032,
				overflow => add_overflow_s032
				);

	Adder_Signed_20bits_033 : Adder_Signed_20bits
	port map(	input_a => multi_s66,
				input_b => multi_s67,
				output => add_output_s033,
				overflow => add_overflow_s033
				);

	Adder_Signed_20bits_034 : Adder_Signed_20bits
	port map(	input_a => multi_s68,
				input_b => multi_s69,
				output => add_output_s034,
				overflow => add_overflow_s034
				);

	Adder_Signed_20bits_035 : Adder_Signed_20bits
	port map(	input_a => multi_s70,
				input_b => b,
				output => add_output_s035,
				overflow => add_overflow_s035
				);

	Adder_Signed_20bits_10 : Adder_Signed_20bits
	port map(	input_a => add_output_s00,
				input_b => add_output_s01,
				output => add_output_s10,
				overflow => add_overflow_s10
				);

	Adder_Signed_20bits_11 : Adder_Signed_20bits
	port map(	input_a => add_output_s02,
				input_b => add_output_s03,
				output => add_output_s11,
				overflow => add_overflow_s11
				);

	Adder_Signed_20bits_12 : Adder_Signed_20bits
	port map(	input_a => add_output_s04,
				input_b => add_output_s05,
				output => add_output_s12,
				overflow => add_overflow_s12
				);

	Adder_Signed_20bits_13 : Adder_Signed_20bits
	port map(	input_a => add_output_s06,
				input_b => add_output_s07,
				output => add_output_s13,
				overflow => add_overflow_s13
				);

	Adder_Signed_20bits_14 : Adder_Signed_20bits
	port map(	input_a => add_output_s08,
				input_b => add_output_s09,
				output => add_output_s14,
				overflow => add_overflow_s14
				);

	Adder_Signed_20bits_15 : Adder_Signed_20bits
	port map(	input_a => add_output_s010,
				input_b => add_output_s011,
				output => add_output_s15,
				overflow => add_overflow_s15
				);

	Adder_Signed_20bits_16 : Adder_Signed_20bits
	port map(	input_a => add_output_s012,
				input_b => add_output_s013,
				output => add_output_s16,
				overflow => add_overflow_s16
				);

	Adder_Signed_20bits_17 : Adder_Signed_20bits
	port map(	input_a => add_output_s014,
				input_b => add_output_s015,
				output => add_output_s17,
				overflow => add_overflow_s17
				);

	Adder_Signed_20bits_18 : Adder_Signed_20bits
	port map(	input_a => add_output_s016,
				input_b => add_output_s017,
				output => add_output_s18,
				overflow => add_overflow_s18
				);

	Adder_Signed_20bits_19 : Adder_Signed_20bits
	port map(	input_a => add_output_s018,
				input_b => add_output_s019,
				output => add_output_s19,
				overflow => add_overflow_s19
				);

	Adder_Signed_20bits_110 : Adder_Signed_20bits
	port map(	input_a => add_output_s020,
				input_b => add_output_s021,
				output => add_output_s110,
				overflow => add_overflow_s110
				);

	Adder_Signed_20bits_111 : Adder_Signed_20bits
	port map(	input_a => add_output_s022,
				input_b => add_output_s023,
				output => add_output_s111,
				overflow => add_overflow_s111
				);

	Adder_Signed_20bits_112 : Adder_Signed_20bits
	port map(	input_a => add_output_s024,
				input_b => add_output_s025,
				output => add_output_s112,
				overflow => add_overflow_s112
				);

	Adder_Signed_20bits_113 : Adder_Signed_20bits
	port map(	input_a => add_output_s026,
				input_b => add_output_s027,
				output => add_output_s113,
				overflow => add_overflow_s113
				);

	Adder_Signed_20bits_114 : Adder_Signed_20bits
	port map(	input_a => add_output_s028,
				input_b => add_output_s029,
				output => add_output_s114,
				overflow => add_overflow_s114
				);

	Adder_Signed_20bits_115 : Adder_Signed_20bits
	port map(	input_a => add_output_s030,
				input_b => add_output_s031,
				output => add_output_s115,
				overflow => add_overflow_s115
				);

	Adder_Signed_20bits_116 : Adder_Signed_20bits
	port map(	input_a => add_output_s032,
				input_b => add_output_s033,
				output => add_output_s116,
				overflow => add_overflow_s116
				);

	Adder_Signed_20bits_117 : Adder_Signed_20bits
	port map(	input_a => add_output_s034,
				input_b => add_output_s035,
				output => add_output_s117,
				overflow => add_overflow_s117
				);

	Adder_Signed_20bits_20 : Adder_Signed_20bits
	port map(	input_a => add_output_s10,
				input_b => add_output_s11,
				output => add_output_s20,
				overflow => add_overflow_s20
				);

	Adder_Signed_20bits_21 : Adder_Signed_20bits
	port map(	input_a => add_output_s12,
				input_b => add_output_s13,
				output => add_output_s21,
				overflow => add_overflow_s21
				);

	Adder_Signed_20bits_22 : Adder_Signed_20bits
	port map(	input_a => add_output_s14,
				input_b => add_output_s15,
				output => add_output_s22,
				overflow => add_overflow_s22
				);

	Adder_Signed_20bits_23 : Adder_Signed_20bits
	port map(	input_a => add_output_s16,
				input_b => add_output_s17,
				output => add_output_s23,
				overflow => add_overflow_s23
				);

	Adder_Signed_20bits_24 : Adder_Signed_20bits
	port map(	input_a => add_output_s18,
				input_b => add_output_s19,
				output => add_output_s24,
				overflow => add_overflow_s24
				);

	Adder_Signed_20bits_25 : Adder_Signed_20bits
	port map(	input_a => add_output_s110,
				input_b => add_output_s111,
				output => add_output_s25,
				overflow => add_overflow_s25
				);

	Adder_Signed_20bits_26 : Adder_Signed_20bits
	port map(	input_a => add_output_s112,
				input_b => add_output_s113,
				output => add_output_s26,
				overflow => add_overflow_s26
				);

	Adder_Signed_20bits_27 : Adder_Signed_20bits
	port map(	input_a => add_output_s114,
				input_b => add_output_s115,
				output => add_output_s27,
				overflow => add_overflow_s27
				);

	Adder_Signed_20bits_28 : Adder_Signed_20bits
	port map(	input_a => add_output_s116,
				input_b => add_output_s117,
				output => add_output_s28,
				overflow => add_overflow_s28
				);

	Adder_Signed_20bits_30 : Adder_Signed_20bits
	port map(	input_a => add_output_s20,
				input_b => add_output_s21,
				output => add_output_s30,
				overflow => add_overflow_s30
				);

	Adder_Signed_20bits_31 : Adder_Signed_20bits
	port map(	input_a => add_output_s22,
				input_b => add_output_s23,
				output => add_output_s31,
				overflow => add_overflow_s31
				);

	Adder_Signed_20bits_32 : Adder_Signed_20bits
	port map(	input_a => add_output_s24,
				input_b => add_output_s25,
				output => add_output_s32,
				overflow => add_overflow_s32
				);

	Adder_Signed_20bits_33 : Adder_Signed_20bits
	port map(	input_a => add_output_s26,
				input_b => add_output_s27,
				output => add_output_s33,
				overflow => add_overflow_s33
				);

	Adder_Signed_20bits_40 : Adder_Signed_20bits
	port map(	input_a => add_output_s30,
				input_b => add_output_s31,
				output => add_output_s40,
				overflow => add_overflow_s40
				);

	Adder_Signed_20bits_41 : Adder_Signed_20bits
	port map(	input_a => add_output_s32,
				input_b => add_output_s33,
				output => add_output_s41,
				overflow => add_overflow_s41
				);

	Adder_Signed_20bits_50 : Adder_Signed_20bits
	port map(	input_a => add_output_s40,
				input_b => add_output_s41,
				output => add_output_s50,
				overflow => add_overflow_s50
				);

	Adder_Signed_20bits_60 : Adder_Signed_20bits
	port map(	input_a => add_output_s50,
				input_b => add_output_s28,
				output => add_output_s60,
				overflow => add_overflow_s60
				);






end Behavioral;